// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Fri May  8 21:56:50 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [7:0] LEGUP_0 = 8'd0;
parameter [7:0] LEGUP_F_main_BB_entry_1 = 8'd1;
parameter [7:0] LEGUP_F_main_BB_entry_2 = 8'd2;
parameter [7:0] LEGUP_F_main_BB_entry_3 = 8'd3;
parameter [7:0] LEGUP_F_main_BB_entry_4 = 8'd4;
parameter [7:0] LEGUP_F_main_BB_entry_5 = 8'd5;
parameter [7:0] LEGUP_F_main_BB_entry_6 = 8'd6;
parameter [7:0] LEGUP_F_main_BB_entry_7 = 8'd7;
parameter [7:0] LEGUP_F_main_BB_entry_8 = 8'd8;
parameter [7:0] LEGUP_F_main_BB_entry_9 = 8'd9;
parameter [7:0] LEGUP_F_main_BB_entry_10 = 8'd10;
parameter [7:0] LEGUP_F_main_BB_entry_11 = 8'd11;
parameter [7:0] LEGUP_F_main_BB_entry_12 = 8'd12;
parameter [7:0] LEGUP_F_main_BB_entry_13 = 8'd13;
parameter [7:0] LEGUP_F_main_BB_entry_14 = 8'd14;
parameter [7:0] LEGUP_F_main_BB_entry_15 = 8'd15;
parameter [7:0] LEGUP_F_main_BB_entry_16 = 8'd16;
parameter [7:0] LEGUP_F_main_BB_entry_17 = 8'd17;
parameter [7:0] LEGUP_F_main_BB_entry_18 = 8'd18;
parameter [7:0] LEGUP_F_main_BB_entry_19 = 8'd19;
parameter [7:0] LEGUP_F_main_BB_entry_20 = 8'd20;
parameter [7:0] LEGUP_F_main_BB_entry_21 = 8'd21;
parameter [7:0] LEGUP_F_main_BB_entry_22 = 8'd22;
parameter [7:0] LEGUP_F_main_BB_entry_23 = 8'd23;
parameter [7:0] LEGUP_F_main_BB_entry_24 = 8'd24;
parameter [7:0] LEGUP_F_main_BB_entry_25 = 8'd25;
parameter [7:0] LEGUP_F_main_BB_entry_26 = 8'd26;
parameter [7:0] LEGUP_F_main_BB_entry_27 = 8'd27;
parameter [7:0] LEGUP_F_main_BB_entry_28 = 8'd28;
parameter [7:0] LEGUP_F_main_BB_entry_29 = 8'd29;
parameter [7:0] LEGUP_F_main_BB_entry_30 = 8'd30;
parameter [7:0] LEGUP_F_main_BB_entry_31 = 8'd31;
parameter [7:0] LEGUP_F_main_BB_entry_32 = 8'd32;
parameter [7:0] LEGUP_F_main_BB_entry_33 = 8'd33;
parameter [7:0] LEGUP_F_main_BB_entry_34 = 8'd34;
parameter [7:0] LEGUP_F_main_BB_entry_35 = 8'd35;
parameter [7:0] LEGUP_F_main_BB_entry_36 = 8'd36;
parameter [7:0] LEGUP_F_main_BB_entry_37 = 8'd37;
parameter [7:0] LEGUP_F_main_BB_entry_38 = 8'd38;
parameter [7:0] LEGUP_F_main_BB_entry_39 = 8'd39;
parameter [7:0] LEGUP_F_main_BB_entry_40 = 8'd40;
parameter [7:0] LEGUP_F_main_BB_entry_41 = 8'd41;
parameter [7:0] LEGUP_F_main_BB_entry_42 = 8'd42;
parameter [7:0] LEGUP_F_main_BB_entry_43 = 8'd43;
parameter [7:0] LEGUP_F_main_BB_for_cond171_preheader_44 = 8'd44;
parameter [7:0] LEGUP_F_main_BB_for_cond171_preheader_45 = 8'd45;
parameter [7:0] LEGUP_F_main_BB_for_body173_46 = 8'd46;
parameter [7:0] LEGUP_F_main_BB_for_body173_47 = 8'd47;
parameter [7:0] LEGUP_F_main_BB_if_then_48 = 8'd48;
parameter [7:0] LEGUP_F_main_BB_if_then_49 = 8'd49;
parameter [7:0] LEGUP_F_main_BB_for_inc_50 = 8'd50;
parameter [7:0] LEGUP_F_main_BB_for_inc178_51 = 8'd51;
parameter [7:0] LEGUP_F_main_BB_for_cond186_preheader_preheader_52 = 8'd52;
parameter [7:0] LEGUP_F_main_BB_for_cond186_preheader_53 = 8'd53;
parameter [7:0] LEGUP_F_main_BB_for_cond186_preheader_54 = 8'd54;
parameter [7:0] LEGUP_F_main_BB_for_body188_55 = 8'd55;
parameter [7:0] LEGUP_F_main_BB_for_body188_56 = 8'd56;
parameter [7:0] LEGUP_F_main_BB_if_then192_57 = 8'd57;
parameter [7:0] LEGUP_F_main_BB_if_then192_58 = 8'd58;
parameter [7:0] LEGUP_F_main_BB_for_inc195_59 = 8'd59;
parameter [7:0] LEGUP_F_main_BB_for_inc198_60 = 8'd60;
parameter [7:0] LEGUP_F_main_BB_for_body203_preheader_61 = 8'd61;
parameter [7:0] LEGUP_F_main_BB_for_body203_62 = 8'd62;
parameter [7:0] LEGUP_F_main_BB_for_body203_63 = 8'd63;
parameter [7:0] LEGUP_F_main_BB_for_body208_64 = 8'd64;
parameter [7:0] LEGUP_F_main_BB_for_body208_65 = 8'd65;
parameter [7:0] LEGUP_F_main_BB_for_inc214_66 = 8'd66;
parameter [7:0] LEGUP_F_main_BB_for_cond220_preheader_preheader_67 = 8'd67;
parameter [7:0] LEGUP_F_main_BB_for_cond220_preheader_68 = 8'd68;
parameter [7:0] LEGUP_F_main_BB_for_cond220_preheader_69 = 8'd69;
parameter [7:0] LEGUP_F_main_BB_for_body222_us_preheader_70 = 8'd70;
parameter [7:0] LEGUP_F_main_BB_for_body222_us_71 = 8'd71;
parameter [7:0] LEGUP_F_main_BB_for_body222_us_72 = 8'd72;
parameter [7:0] LEGUP_F_main_BB_for_body222_us_73 = 8'd73;
parameter [7:0] LEGUP_F_main_BB_if_then226_us_74 = 8'd74;
parameter [7:0] LEGUP_F_main_BB_if_then226_us_75 = 8'd75;
parameter [7:0] LEGUP_F_main_BB_if_then226_us_76 = 8'd76;
parameter [7:0] LEGUP_F_main_BB_if_then226_us_77 = 8'd77;
parameter [7:0] LEGUP_F_main_BB_for_inc291_us_78 = 8'd78;
parameter [7:0] LEGUP_F_main_BB_for_inc291_us_79 = 8'd79;
parameter [7:0] LEGUP_F_main_BB_for_inc291_us_80 = 8'd80;
parameter [7:0] LEGUP_F_main_BB_for_inc294_loopexit_81 = 8'd81;
parameter [7:0] LEGUP_F_main_BB_for_inc294_82 = 8'd82;
parameter [7:0] LEGUP_F_main_BB_for_body300_preheader_83 = 8'd83;
parameter [7:0] LEGUP_F_main_BB_for_body300_84 = 8'd84;
parameter [7:0] LEGUP_F_main_BB_for_body300_85 = 8'd85;
parameter [7:0] LEGUP_F_main_BB_for_body_i_86 = 8'd86;
parameter [7:0] LEGUP_F_main_BB_for_body_i_87 = 8'd87;
parameter [7:0] LEGUP_F_main_BB_for_end_i_88 = 8'd88;
parameter [7:0] LEGUP_F_main_BB_for_end_i_89 = 8'd89;
parameter [7:0] LEGUP_F_main_BB_for_body6_i_90 = 8'd90;
parameter [7:0] LEGUP_F_main_BB_for_body_i_i_91 = 8'd91;
parameter [7:0] LEGUP_F_main_BB_for_body_i_i_92 = 8'd92;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true_i_i_93 = 8'd93;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true_i_i_94 = 8'd94;
parameter [7:0] LEGUP_F_main_BB_for_inc_i_i_95 = 8'd95;
parameter [7:0] LEGUP_F_main_BB_minDistance_exit_i_96 = 8'd96;
parameter [7:0] LEGUP_F_main_BB_minDistance_exit_i_97 = 8'd97;
parameter [7:0] LEGUP_F_main_BB_for_body11_i_98 = 8'd98;
parameter [7:0] LEGUP_F_main_BB_for_body11_i_99 = 8'd99;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true_i_100 = 8'd100;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true_i_101 = 8'd101;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true16_i_102 = 8'd102;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true16_i_103 = 8'd103;
parameter [7:0] LEGUP_F_main_BB_if_then_i_104 = 8'd104;
parameter [7:0] LEGUP_F_main_BB_if_then_i_105 = 8'd105;
parameter [7:0] LEGUP_F_main_BB_for_inc28_i_106 = 8'd106;
parameter [7:0] LEGUP_F_main_BB_for_inc31_i_107 = 8'd107;
parameter [7:0] LEGUP_F_main_BB_dijkstra_exit_108 = 8'd108;
parameter [7:0] LEGUP_F_main_BB_dijkstra_exit_109 = 8'd109;
parameter [7:0] LEGUP_F_main_BB_if_end313_preheader_110 = 8'd110;
parameter [7:0] LEGUP_F_main_BB_if_end313_111 = 8'd111;
parameter [7:0] LEGUP_F_main_BB_if_end313_112 = 8'd112;
parameter [7:0] LEGUP_F_main_BB_if_then322_113 = 8'd113;
parameter [7:0] LEGUP_F_main_BB_if_then322_114 = 8'd114;
parameter [7:0] LEGUP_F_main_BB_for_inc340_loopexit_115 = 8'd115;
parameter [7:0] LEGUP_F_main_BB_for_inc340_116 = 8'd116;
parameter [7:0] LEGUP_F_main_BB_for_end342_loopexit_117 = 8'd117;
parameter [7:0] LEGUP_F_main_BB_for_end342_loopexit1_118 = 8'd118;
parameter [7:0] LEGUP_F_main_BB_for_end342_119 = 8'd119;
parameter [7:0] LEGUP_F_main_BB_for_inc291_8_120 = 8'd120;
parameter [7:0] LEGUP_F_main_BB_for_inc291_8_121 = 8'd121;
parameter [7:0] LEGUP_F_main_BB_for_inc291_8_122 = 8'd122;
parameter [7:0] LEGUP_F_main_BB_for_inc291_8_123 = 8'd123;
parameter [7:0] LEGUP_F_main_BB_for_inc291_8_124 = 8'd124;
parameter [7:0] LEGUP_F_main_BB_for_inc291_8_125 = 8'd125;
parameter [7:0] LEGUP_F_main_BB_for_inc291_8_126 = 8'd126;
parameter [7:0] LEGUP_F_main_BB_for_inc291_8_127 = 8'd127;
parameter [7:0] LEGUP_F_main_BB_for_inc291_8_128 = 8'd128;
parameter [7:0] LEGUP_F_main_BB_for_inc291_8_129 = 8'd129;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [7:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [7:0] next_state;
wire  fsm_stall;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_vla1422_sub;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_vla421_sub;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx3;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx4;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx5_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx6_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx7;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx7_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx8;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx8_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx9;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx9_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx10;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx10_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx11;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx11_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx12;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx12_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx13;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx13_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx14;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx14_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx15;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx15_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx16;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx16_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx17;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx17_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx18;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx18_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx19;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx19_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx20;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx20_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx21;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx21_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx22;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx22_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx23;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx23_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx24;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx24_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx25;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx25_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx26;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx26_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx27;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx27_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx28;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx28_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx29;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx29_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx30;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx30_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx31;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx31_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx32;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx32_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx33;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx33_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx34;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx34_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx35;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx35_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx36;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx36_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx37;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx37_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx38;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx38_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx39;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx39_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx40;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx40_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx41;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx41_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx42;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx42_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx43;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx43_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx44;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx44_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx45;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx45_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx46;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx46_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx47;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx47_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx48;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx48_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx49;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx49_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx50;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx50_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx51;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx51_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx52;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx52_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx53;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx53_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx54;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx54_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx55;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx55_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx56;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx56_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx57;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx57_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx58;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx58_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx59;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx59_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx60;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx60_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx61;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx61_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx62;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx62_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx63;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx63_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx64;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx64_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx65;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx65_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx66;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx66_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx67;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx67_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx68;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx68_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx69;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx69_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx70;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx70_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx71;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx71_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx72;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx72_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx73;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx73_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx74;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx74_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx75;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx75_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx76;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx76_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx77;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx77_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx78;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx78_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx79;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx79_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx80;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx80_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx81;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx81_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx82;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx82_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx83;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx83_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx84;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx84_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx85;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx85_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx86;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx86_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx87;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx87_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx88;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx88_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx89;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx89_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx90;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx90_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx91;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx91_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx92;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx92_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx93;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx93_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx94;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx94_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx95;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx95_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx96;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx96_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx97;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx97_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx98;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx98_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx99;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx99_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx100;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx100_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx101;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx101_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx102;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx102_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx103;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx103_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx104;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx104_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx105;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx105_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx106;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx106_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx107;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx107_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx108;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx108_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx109;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx109_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx110;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx110_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx111;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx111_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx112;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx112_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx113;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx113_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx114;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx114_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx115;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx115_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx116;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx116_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx117;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx117_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx118;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx118_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx119;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx119_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx120;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx120_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx121;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx121_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx122;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx122_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx123;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx123_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx124;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx124_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx125;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx125_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx126;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx126_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx127;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx127_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx128;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx128_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx129;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx129_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx130;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx130_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx131;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx131_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx132;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx132_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx133;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx133_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx134;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx134_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx135;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx135_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx136;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx136_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx137;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx137_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx138;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx138_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx139;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx139_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx140;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx140_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx141;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx141_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx142;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx142_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx143;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx143_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx144;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx144_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx145;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx145_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx146;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx146_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx147;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx147_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx148;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx148_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx149;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx149_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx150;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx150_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx151;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx151_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx152;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx152_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx153;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx153_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx154;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx154_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx155;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx155_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx156;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx156_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx157;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx157_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx158;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx158_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx159;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx159_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx160;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx160_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx161;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx161_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx162;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx162_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx163;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx163_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx164;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx164_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx165;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx165_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx166;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx166_reg;
reg [6:0] main_for_cond171_preheader_j169_0444;
reg [6:0] main_for_cond171_preheader_j169_0444_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond171_preheader_arrayidx174;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond171_preheader_arrayidx177;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond171_preheader_arrayidx177_reg;
reg [31:0] main_for_cond171_preheader_0;
reg [31:0] main_for_cond171_preheader_0_reg;
reg [31:0] main_for_body173_1;
reg [31:0] main_for_body173_1_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body173_arrayidx175;
reg [31:0] main_for_body173_2;
reg  main_for_body173_cmp176;
reg [31:0] main_for_inc_3;
reg  main_for_inc_exitcond11;
reg [7:0] main_for_inc178_4;
reg  main_for_inc178_exitcond12;
reg [6:0] main_for_cond186_preheader_j181_0442;
reg [6:0] main_for_cond186_preheader_j181_0442_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond186_preheader_arrayidx189;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond186_preheader_arrayidx193;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond186_preheader_arrayidx193_reg;
reg [31:0] main_for_cond186_preheader_5;
reg [31:0] main_for_cond186_preheader_5_reg;
reg [31:0] main_for_body188_6;
reg [31:0] main_for_body188_6_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body188_arrayidx190;
reg [31:0] main_for_body188_7;
reg  main_for_body188_cmp191;
reg [31:0] main_for_inc195_8;
reg  main_for_inc195_exitcond;
reg [7:0] main_for_inc198_9;
reg  main_for_inc198_exitcond10;
reg [6:0] main_for_body203_i_0440;
reg [6:0] main_for_body203_i_0440_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body203_arrayidx204;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body203_arrayidx205;
reg [31:0] main_for_body208_j_0439;
reg [31:0] main_for_body208_j_0439_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body208_arrayidx210;
reg [31:0] main_for_body208_10;
reg [31:0] main_for_body208_10_reg;
reg  main_for_body208_exitcond8;
reg  main_for_body208_exitcond8_reg;
reg [7:0] main_for_inc214_11;
reg  main_for_inc214_exitcond9;
reg [3:0] main_for_cond220_preheader_12;
reg [3:0] main_for_cond220_preheader_12_reg;
reg [30:0] main_for_cond220_preheader_bit_select13;
reg [23:0] main_for_cond220_preheader_bit_select9;
reg [22:0] main_for_cond220_preheader_bit_select7;
reg [4:0] main_for_cond220_preheader_sr_negate;
reg [26:0] main_for_cond220_preheader_bit_select11;
reg [31:0] main_for_cond220_preheader_bit_concat14;
reg [31:0] main_for_cond220_preheader_bit_concat12;
reg [31:0] main_for_cond220_preheader_bit_concat10;
reg [31:0] main_for_cond220_preheader_bit_concat8;
reg [31:0] main_for_cond220_preheader_sr_add;
reg [31:0] main_for_cond220_preheader_sr_add_reg;
reg [31:0] main_for_cond220_preheader_sr_add16;
reg [31:0] main_for_cond220_preheader_sr_add16_reg;
reg [31:0] main_for_cond220_preheader_sr_add17;
reg [31:0] main_for_cond220_preheader_sr_add17_reg;
reg [30:0] main_for_cond220_preheader_bit_select5;
reg [31:0] main_for_cond220_preheader_13;
reg [31:0] main_for_cond220_preheader_13_reg;
reg [31:0] main_for_cond220_preheader_bit_concat6;
reg [31:0] main_for_cond220_preheader_bit_concat6_reg;
reg [31:0] main_for_cond220_preheader_14;
reg [31:0] main_for_cond220_preheader_14_reg;
reg [31:0] main_for_cond220_preheader_15;
reg [31:0] main_for_cond220_preheader_15_reg;
reg [31:0] main_for_cond220_preheader_16;
reg [31:0] main_for_cond220_preheader_16_reg;
reg [31:0] main_for_cond220_preheader_17;
reg [31:0] main_for_cond220_preheader_17_reg;
reg [31:0] main_for_cond220_preheader_18;
reg [31:0] main_for_cond220_preheader_18_reg;
reg [31:0] main_for_cond220_preheader_19;
reg [31:0] main_for_cond220_preheader_19_reg;
reg  main_for_cond220_preheader_cmp223;
reg  main_for_cond220_preheader_cmp223_reg;
reg [31:0] main_for_body222_us_20;
reg [31:0] main_for_body222_us_20_reg;
reg [30:0] main_for_body222_us_bit_select3;
reg [27:0] main_for_body222_us_bit_select1;
reg [25:0] main_for_body222_us_bit_select;
reg [31:0] main_for_body222_us_bit_concat4;
reg [31:0] main_for_body222_us_bit_concat2;
reg [31:0] main_for_body222_us_bit_concat;
reg [31:0] main_for_body222_us_sr_add21;
reg [31:0] main_for_body222_us_sr_add22;
reg [31:0] main_for_body222_us_sr_add22_reg;
reg [31:0] main_for_body222_us_21;
reg [31:0] main_for_body222_us_21_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body222_us_arrayidx262_us;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body222_us_arrayidx262_us_reg;
reg [31:0] main_for_body222_us_22;
reg [31:0] main_for_body222_us_22_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body222_us_arrayidx269_us;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body222_us_arrayidx269_us_reg;
reg  main_for_body222_us_cmp224_us;
reg  main_for_body222_us_cmp224_us_reg;
reg [31:0] main_if_then226_us_23;
reg [31:0] main_if_then226_us_23_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then226_us_arrayidx231_us;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then226_us_arrayidx238_us;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then226_us_arrayidx238_us_reg;
reg [31:0] main_for_inc291_us_24;
reg [31:0] main_for_inc291_us_24_reg;
reg  main_for_inc291_us_exitcond6;
reg  main_for_inc291_us_exitcond6_reg;
reg [4:0] main_for_inc294_25;
reg  main_for_inc294_exitcond7;
reg [6:0] main_for_body300_i_2435;
reg [6:0] main_for_body300_i_2435_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body300_arrayidx301;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body300_arrayidx302;
reg [7:0] main_for_body300_inc341;
reg [7:0] main_for_body300_inc341_reg;
reg [31:0] main_for_body300_26;
reg [31:0] main_for_body300_26_reg;
reg [31:0] main_for_body300_27;
reg [31:0] main_for_body300_27_reg;
reg [31:0] main_for_body_i_i_057_i;
reg [31:0] main_for_body_i_i_057_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx1_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx2_i;
reg [31:0] main_for_body_i_28;
reg [31:0] main_for_body_i_28_reg;
reg  main_for_body_i_exitcond2;
reg  main_for_body_i_exitcond2_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_end_i_arrayidx_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_end_i_arrayidx3_i;
reg [31:0] main_for_body6_i_count_056_i;
reg [31:0] main_for_body6_i_count_056_i_reg;
reg [31:0] main_for_body_i_i_29;
reg [31:0] main_for_body_i_i_29_reg;
reg [31:0] main_for_body_i_i_min_index_012_i_i;
reg [31:0] main_for_body_i_i_min_index_012_i_i_reg;
reg [31:0] main_for_body_i_i_min_011_i_i;
reg [31:0] main_for_body_i_i_min_011_i_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_i_arrayidx_i_i;
reg [31:0] main_for_body_i_i_30;
reg  main_for_body_i_i_cmp1_i_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_land_lhs_true_i_i_arrayidx2_i_i;
reg [31:0] main_land_lhs_true_i_i_31;
reg  main_land_lhs_true_i_i_cmp3_i_i;
reg [31:0] main_land_lhs_true_i_i_min_0_i_i;
reg [31:0] main_land_lhs_true_i_i_min_index_0_v_0_i_i;
reg [31:0] main_for_inc_i_i_min_1_i_i;
reg [31:0] main_for_inc_i_i_min_1_i_i_reg;
reg [31:0] main_for_inc_i_i_min_index_1_i_i;
reg [31:0] main_for_inc_i_i_min_index_1_i_i_reg;
reg [31:0] main_for_inc_i_i_32;
reg  main_for_inc_i_i_exitcond3;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_minDistance_exit_i_arrayidx8_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_minDistance_exit_i_arrayidx17_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_minDistance_exit_i_arrayidx17_i_reg;
reg [31:0] main_for_body11_i_v_055_i;
reg [31:0] main_for_body11_i_v_055_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx12_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx20_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx20_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx22_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx22_i_reg;
reg [31:0] main_for_body11_i_33;
reg  main_for_body11_i_tobool_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_land_lhs_true_i_arrayidx14_i;
reg [31:0] main_land_lhs_true_i_34;
reg [31:0] main_land_lhs_true_i_34_reg;
reg  main_land_lhs_true_i_tobool15_i;
reg [31:0] main_land_lhs_true16_i_35;
reg [31:0] main_land_lhs_true16_i_add_i;
reg [31:0] main_land_lhs_true16_i_add_i_reg;
reg [31:0] main_land_lhs_true16_i_36;
reg  main_land_lhs_true16_i_cmp21_i;
reg [31:0] main_for_inc28_i_37;
reg  main_for_inc28_i_exitcond4;
reg [31:0] main_for_inc31_i_38;
reg  main_for_inc31_i_exitcond5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_dijkstra_exit_arrayidx309431;
reg [31:0] main_dijkstra_exit_39;
reg [31:0] main_dijkstra_exit_39_reg;
reg  main_dijkstra_exit_cmp310432;
reg [31:0] main_if_end313_40;
reg [31:0] main_if_end313_40_reg;
reg [31:0] main_if_end313_origem_1434;
reg [31:0] main_if_end313_origem_1434_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end313_arrayidx314;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end313_arrayidx314_reg;
reg [31:0] main_if_end313_41;
reg [31:0] main_if_end313_41_reg;
reg  main_if_end313_cmp315;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end313_arrayidx317;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end313_arrayidx317_reg;
reg [31:0] main_if_end313_42;
reg [31:0] main_if_end313_42_reg;
reg  main_if_end313_cmp318;
reg  main_if_end313_and320425;
reg [31:0] main_if_then322_add330;
reg [31:0] main_if_then322_add332;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then322_arrayidx309;
reg [31:0] main_if_then322_43;
reg  main_if_then322_cmp310;
reg  main_for_inc340_cmp298;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_1;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_1_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_7;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_7_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_6_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_6_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_5_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_5_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_4_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_4_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_3;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_3_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_3;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_3_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_2;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_2_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_2;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx287_2_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_1;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_1_reg;
reg [31:0] main_for_inc291_8_44;
reg [31:0] main_for_inc291_8_44_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_7;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc291_8_arrayidx280_7_reg;
reg [6:0] main_grid_address_a;
wire [31:0] main_grid_out_a;
wire [6:0] main_grid_address_b;
wire [31:0] main_grid_out_b;
reg [6:0] main_entry_dist_i_address_a;
reg  main_entry_dist_i_write_enable_a;
reg [31:0] main_entry_dist_i_in_a;
wire [31:0] main_entry_dist_i_out_a;
reg [6:0] main_entry_dist_i_address_b;
reg  main_entry_dist_i_write_enable_b;
reg [31:0] main_entry_dist_i_in_b;
wire [31:0] main_entry_dist_i_out_b;
reg [6:0] main_entry_sptSet_i_address_a;
reg  main_entry_sptSet_i_write_enable_a;
reg [31:0] main_entry_sptSet_i_in_a;
wire [31:0] main_entry_sptSet_i_out_a;
reg [6:0] main_entry_parent_address_a;
reg  main_entry_parent_write_enable_a;
reg [31:0] main_entry_parent_in_a;
wire [31:0] main_entry_parent_out_a;
reg [12:0] main_entry_m_address_a;
reg  main_entry_m_write_enable_a;
reg [31:0] main_entry_m_in_a;
wire [31:0] main_entry_m_out_a;
reg [12:0] main_entry_m_address_b;
reg  main_entry_m_write_enable_b;
reg [31:0] main_entry_m_in_b;
wire [31:0] main_entry_m_out_b;
reg [6:0] main_entry_indice_e_address_a;
reg  main_entry_indice_e_write_enable_a;
reg [31:0] main_entry_indice_e_in_a;
wire [31:0] main_entry_indice_e_out_a;
reg [6:0] main_entry_indice_s_address_a;
reg  main_entry_indice_s_write_enable_a;
reg [31:0] main_entry_indice_s_in_a;
wire [31:0] main_entry_indice_s_out_a;
reg [6:0] main_entry_vla421_address_a;
reg  main_entry_vla421_write_enable_a;
reg [31:0] main_entry_vla421_in_a;
wire [31:0] main_entry_vla421_out_a;
reg [6:0] main_entry_vla421_address_b;
reg  main_entry_vla421_write_enable_b;
reg [31:0] main_entry_vla421_in_b;
wire [31:0] main_entry_vla421_out_b;
reg [6:0] main_entry_vla1422_address_a;
reg  main_entry_vla1422_write_enable_a;
reg [31:0] main_entry_vla1422_in_a;
wire [31:0] main_entry_vla1422_out_a;
reg [6:0] main_entry_vla1422_address_b;
reg  main_entry_vla1422_write_enable_b;
reg [31:0] main_entry_vla1422_in_b;
wire [31:0] main_entry_vla1422_out_b;
reg [6:0] main_entry_vla167423_address_a;
reg  main_entry_vla167423_write_enable_a;
reg [31:0] main_entry_vla167423_in_a;
wire [31:0] main_entry_vla167423_out_a;
reg [6:0] main_entry_vla168424_address_a;
reg  main_entry_vla168424_write_enable_a;
reg [31:0] main_entry_vla168424_in_a;
wire [31:0] main_entry_vla168424_out_a;
reg [30:0] main_for_cond220_preheader_12_reg_width_extended;
reg [26:0] main_for_cond220_preheader_sr_negate_width_extended;
wire  main_for_cond220_preheader_bit_concat14_bit_select_operand_2;
wire [4:0] main_for_cond220_preheader_bit_concat12_bit_select_operand_2;
wire [7:0] main_for_cond220_preheader_bit_concat10_bit_select_operand_2;
wire [8:0] main_for_cond220_preheader_bit_concat8_bit_select_operand_2;
reg [4:0] main_for_cond220_preheader_cmp223_op0_temp;
wire [5:0] main_for_cond220_preheader_cmp223_op1_temp;
wire  main_for_cond220_preheader_bit_concat6_bit_select_operand_2;
wire  main_for_body222_us_bit_concat4_bit_select_operand_2;
wire [3:0] main_for_body222_us_bit_concat2_bit_select_operand_2;
wire [5:0] main_for_body222_us_bit_concat_bit_select_operand_2;
wire [5:0] main_for_body222_us_cmp224_us_op1_temp;
wire [4:0] main_if_end313_cmp315_op1_temp;
wire [4:0] main_if_end313_cmp318_op1_temp;
reg [8:0] main_for_inc340_cmp298_op0_temp;
wire [8:0] main_for_inc340_cmp298_op1_temp;



// @main.grid = private unnamed_addr constant [81 x i32] [i32 255, i32 5, i32 9, i32 21, i32 19, i32 45, i32 18, i32 29, i32 67, i32 255, i32 17, i32 4, i32 32, i32 6, i32 51, i32 38, i32 65, i32 66, i32...
rom_dual_port main_grid (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_grid_address_a ),
	.q_a( main_grid_out_a ),
	.address_b( main_grid_address_b ),
	.q_b( main_grid_out_b )
);
defparam main_grid.width_a = 32;
defparam main_grid.widthad_a = 7;
defparam main_grid.numwords_a = 81;
defparam main_grid.width_b = 32;
defparam main_grid.widthad_b = 7;
defparam main_grid.numwords_b = 81;
defparam main_grid.latency = 1;
defparam main_grid.init_file = {`MEM_INIT_DIR, "main_grid.mif"};


//   %dist.i = alloca [81 x i32], align 4, !dbg !83, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_dist_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_dist_i_address_a ),
	.wren_a( main_entry_dist_i_write_enable_a ),
	.data_a( main_entry_dist_i_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_dist_i_out_a ),
	.address_b( main_entry_dist_i_address_b ),
	.wren_b( main_entry_dist_i_write_enable_b ),
	.data_b( main_entry_dist_i_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_dist_i_out_b )
);
defparam main_entry_dist_i.width_a = 32;
defparam main_entry_dist_i.widthad_a = 7;
defparam main_entry_dist_i.width_be_a = 4;
defparam main_entry_dist_i.numwords_a = 81;
defparam main_entry_dist_i.width_b = 32;
defparam main_entry_dist_i.widthad_b = 7;
defparam main_entry_dist_i.width_be_b = 4;
defparam main_entry_dist_i.numwords_b = 81;
defparam main_entry_dist_i.latency = 1;


//   %sptSet.i = alloca [81 x i32], align 4, !dbg !83, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_sptSet_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_sptSet_i_address_a ),
	.wren_a( main_entry_sptSet_i_write_enable_a ),
	.data_a( main_entry_sptSet_i_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_sptSet_i_out_a )
);
defparam main_entry_sptSet_i.width_a = 32;
defparam main_entry_sptSet_i.widthad_a = 7;
defparam main_entry_sptSet_i.width_be_a = 4;
defparam main_entry_sptSet_i.numwords_a = 81;
defparam main_entry_sptSet_i.latency = 1;


//   %parent = alloca [81 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_parent (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_parent_address_a ),
	.wren_a( main_entry_parent_write_enable_a ),
	.data_a( main_entry_parent_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_parent_out_a )
);
defparam main_entry_parent.width_a = 32;
defparam main_entry_parent.widthad_a = 7;
defparam main_entry_parent.width_be_a = 4;
defparam main_entry_parent.numwords_a = 81;
defparam main_entry_parent.latency = 1;


//   %m = alloca [81 x [81 x i32]], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_m (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_m_address_a ),
	.wren_a( main_entry_m_write_enable_a ),
	.data_a( main_entry_m_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_m_out_a ),
	.address_b( main_entry_m_address_b ),
	.wren_b( main_entry_m_write_enable_b ),
	.data_b( main_entry_m_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_m_out_b )
);
defparam main_entry_m.width_a = 32;
defparam main_entry_m.widthad_a = 13;
defparam main_entry_m.width_be_a = 4;
defparam main_entry_m.numwords_a = 6561;
defparam main_entry_m.width_b = 32;
defparam main_entry_m.widthad_b = 13;
defparam main_entry_m.width_be_b = 4;
defparam main_entry_m.numwords_b = 6561;
defparam main_entry_m.latency = 1;


//   %indice_e = alloca [81 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_indice_e (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_indice_e_address_a ),
	.wren_a( main_entry_indice_e_write_enable_a ),
	.data_a( main_entry_indice_e_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_indice_e_out_a )
);
defparam main_entry_indice_e.width_a = 32;
defparam main_entry_indice_e.widthad_a = 7;
defparam main_entry_indice_e.width_be_a = 4;
defparam main_entry_indice_e.numwords_a = 81;
defparam main_entry_indice_e.latency = 1;


//   %indice_s = alloca [81 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_indice_s (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_indice_s_address_a ),
	.wren_a( main_entry_indice_s_write_enable_a ),
	.data_a( main_entry_indice_s_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_indice_s_out_a )
);
defparam main_entry_indice_s.width_a = 32;
defparam main_entry_indice_s.widthad_a = 7;
defparam main_entry_indice_s.width_be_a = 4;
defparam main_entry_indice_s.numwords_a = 81;
defparam main_entry_indice_s.latency = 1;


//   %vla421 = alloca [83 x i32], align 4, !dbg !88, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_vla421 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla421_address_a ),
	.wren_a( main_entry_vla421_write_enable_a ),
	.data_a( main_entry_vla421_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla421_out_a ),
	.address_b( main_entry_vla421_address_b ),
	.wren_b( main_entry_vla421_write_enable_b ),
	.data_b( main_entry_vla421_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_vla421_out_b )
);
defparam main_entry_vla421.width_a = 32;
defparam main_entry_vla421.widthad_a = 7;
defparam main_entry_vla421.width_be_a = 4;
defparam main_entry_vla421.numwords_a = 83;
defparam main_entry_vla421.width_b = 32;
defparam main_entry_vla421.widthad_b = 7;
defparam main_entry_vla421.width_be_b = 4;
defparam main_entry_vla421.numwords_b = 83;
defparam main_entry_vla421.latency = 1;


//   %vla1422 = alloca [83 x i32], align 4, !dbg !89, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_vla1422 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla1422_address_a ),
	.wren_a( main_entry_vla1422_write_enable_a ),
	.data_a( main_entry_vla1422_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla1422_out_a ),
	.address_b( main_entry_vla1422_address_b ),
	.wren_b( main_entry_vla1422_write_enable_b ),
	.data_b( main_entry_vla1422_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_vla1422_out_b )
);
defparam main_entry_vla1422.width_a = 32;
defparam main_entry_vla1422.widthad_a = 7;
defparam main_entry_vla1422.width_be_a = 4;
defparam main_entry_vla1422.numwords_a = 83;
defparam main_entry_vla1422.width_b = 32;
defparam main_entry_vla1422.widthad_b = 7;
defparam main_entry_vla1422.width_be_b = 4;
defparam main_entry_vla1422.numwords_b = 83;
defparam main_entry_vla1422.latency = 1;


//   %vla167423 = alloca [83 x i32], align 4, !dbg !260, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_vla167423 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla167423_address_a ),
	.wren_a( main_entry_vla167423_write_enable_a ),
	.data_a( main_entry_vla167423_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla167423_out_a )
);
defparam main_entry_vla167423.width_a = 32;
defparam main_entry_vla167423.widthad_a = 7;
defparam main_entry_vla167423.width_be_a = 4;
defparam main_entry_vla167423.numwords_a = 83;
defparam main_entry_vla167423.latency = 1;


//   %vla168424 = alloca [83 x i32], align 4, !dbg !260, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_vla168424 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla168424_address_a ),
	.wren_a( main_entry_vla168424_write_enable_a ),
	.data_a( main_entry_vla168424_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla168424_out_a )
);
defparam main_entry_vla168424.width_a = 32;
defparam main_entry_vla168424.widthad_a = 7;
defparam main_entry_vla168424.width_be_a = 4;
defparam main_entry_vla168424.numwords_a = 83;
defparam main_entry_vla168424.latency = 1;

always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_entry_1;
LEGUP_F_main_BB_dijkstra_exit_108:
		next_state = LEGUP_F_main_BB_dijkstra_exit_109;
LEGUP_F_main_BB_dijkstra_exit_109:
	if ((fsm_stall == 1'd0) && (main_dijkstra_exit_cmp310432 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc340_116;
	else if ((fsm_stall == 1'd0) && (main_dijkstra_exit_cmp310432 == 1'd0))
		next_state = LEGUP_F_main_BB_if_end313_preheader_110;
LEGUP_F_main_BB_entry_1:
		next_state = LEGUP_F_main_BB_entry_2;
LEGUP_F_main_BB_entry_10:
		next_state = LEGUP_F_main_BB_entry_11;
LEGUP_F_main_BB_entry_11:
		next_state = LEGUP_F_main_BB_entry_12;
LEGUP_F_main_BB_entry_12:
		next_state = LEGUP_F_main_BB_entry_13;
LEGUP_F_main_BB_entry_13:
		next_state = LEGUP_F_main_BB_entry_14;
LEGUP_F_main_BB_entry_14:
		next_state = LEGUP_F_main_BB_entry_15;
LEGUP_F_main_BB_entry_15:
		next_state = LEGUP_F_main_BB_entry_16;
LEGUP_F_main_BB_entry_16:
		next_state = LEGUP_F_main_BB_entry_17;
LEGUP_F_main_BB_entry_17:
		next_state = LEGUP_F_main_BB_entry_18;
LEGUP_F_main_BB_entry_18:
		next_state = LEGUP_F_main_BB_entry_19;
LEGUP_F_main_BB_entry_19:
		next_state = LEGUP_F_main_BB_entry_20;
LEGUP_F_main_BB_entry_2:
		next_state = LEGUP_F_main_BB_entry_3;
LEGUP_F_main_BB_entry_20:
		next_state = LEGUP_F_main_BB_entry_21;
LEGUP_F_main_BB_entry_21:
		next_state = LEGUP_F_main_BB_entry_22;
LEGUP_F_main_BB_entry_22:
		next_state = LEGUP_F_main_BB_entry_23;
LEGUP_F_main_BB_entry_23:
		next_state = LEGUP_F_main_BB_entry_24;
LEGUP_F_main_BB_entry_24:
		next_state = LEGUP_F_main_BB_entry_25;
LEGUP_F_main_BB_entry_25:
		next_state = LEGUP_F_main_BB_entry_26;
LEGUP_F_main_BB_entry_26:
		next_state = LEGUP_F_main_BB_entry_27;
LEGUP_F_main_BB_entry_27:
		next_state = LEGUP_F_main_BB_entry_28;
LEGUP_F_main_BB_entry_28:
		next_state = LEGUP_F_main_BB_entry_29;
LEGUP_F_main_BB_entry_29:
		next_state = LEGUP_F_main_BB_entry_30;
LEGUP_F_main_BB_entry_3:
		next_state = LEGUP_F_main_BB_entry_4;
LEGUP_F_main_BB_entry_30:
		next_state = LEGUP_F_main_BB_entry_31;
LEGUP_F_main_BB_entry_31:
		next_state = LEGUP_F_main_BB_entry_32;
LEGUP_F_main_BB_entry_32:
		next_state = LEGUP_F_main_BB_entry_33;
LEGUP_F_main_BB_entry_33:
		next_state = LEGUP_F_main_BB_entry_34;
LEGUP_F_main_BB_entry_34:
		next_state = LEGUP_F_main_BB_entry_35;
LEGUP_F_main_BB_entry_35:
		next_state = LEGUP_F_main_BB_entry_36;
LEGUP_F_main_BB_entry_36:
		next_state = LEGUP_F_main_BB_entry_37;
LEGUP_F_main_BB_entry_37:
		next_state = LEGUP_F_main_BB_entry_38;
LEGUP_F_main_BB_entry_38:
		next_state = LEGUP_F_main_BB_entry_39;
LEGUP_F_main_BB_entry_39:
		next_state = LEGUP_F_main_BB_entry_40;
LEGUP_F_main_BB_entry_4:
		next_state = LEGUP_F_main_BB_entry_5;
LEGUP_F_main_BB_entry_40:
		next_state = LEGUP_F_main_BB_entry_41;
LEGUP_F_main_BB_entry_41:
		next_state = LEGUP_F_main_BB_entry_42;
LEGUP_F_main_BB_entry_42:
		next_state = LEGUP_F_main_BB_entry_43;
LEGUP_F_main_BB_entry_43:
		next_state = LEGUP_F_main_BB_for_cond171_preheader_44;
LEGUP_F_main_BB_entry_5:
		next_state = LEGUP_F_main_BB_entry_6;
LEGUP_F_main_BB_entry_6:
		next_state = LEGUP_F_main_BB_entry_7;
LEGUP_F_main_BB_entry_7:
		next_state = LEGUP_F_main_BB_entry_8;
LEGUP_F_main_BB_entry_8:
		next_state = LEGUP_F_main_BB_entry_9;
LEGUP_F_main_BB_entry_9:
		next_state = LEGUP_F_main_BB_entry_10;
LEGUP_F_main_BB_for_body11_i_98:
		next_state = LEGUP_F_main_BB_for_body11_i_99;
LEGUP_F_main_BB_for_body11_i_99:
	if ((fsm_stall == 1'd0) && (main_for_body11_i_tobool_i == 1'd1))
		next_state = LEGUP_F_main_BB_land_lhs_true_i_100;
	else if ((fsm_stall == 1'd0) && (main_for_body11_i_tobool_i == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc28_i_106;
LEGUP_F_main_BB_for_body173_46:
		next_state = LEGUP_F_main_BB_for_body173_47;
LEGUP_F_main_BB_for_body173_47:
	if ((fsm_stall == 1'd0) && (main_for_body173_cmp176 == 1'd1))
		next_state = LEGUP_F_main_BB_if_then_48;
	else if ((fsm_stall == 1'd0) && (main_for_body173_cmp176 == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc_50;
LEGUP_F_main_BB_for_body188_55:
		next_state = LEGUP_F_main_BB_for_body188_56;
LEGUP_F_main_BB_for_body188_56:
	if ((fsm_stall == 1'd0) && (main_for_body188_cmp191 == 1'd1))
		next_state = LEGUP_F_main_BB_if_then192_57;
	else if ((fsm_stall == 1'd0) && (main_for_body188_cmp191 == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc195_59;
LEGUP_F_main_BB_for_body203_62:
		next_state = LEGUP_F_main_BB_for_body203_63;
LEGUP_F_main_BB_for_body203_63:
		next_state = LEGUP_F_main_BB_for_body208_64;
LEGUP_F_main_BB_for_body203_preheader_61:
		next_state = LEGUP_F_main_BB_for_body203_62;
LEGUP_F_main_BB_for_body208_64:
		next_state = LEGUP_F_main_BB_for_body208_65;
LEGUP_F_main_BB_for_body208_65:
	if ((fsm_stall == 1'd0) && (main_for_body208_exitcond8_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc214_66;
	else if ((fsm_stall == 1'd0) && (main_for_body208_exitcond8_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body208_64;
LEGUP_F_main_BB_for_body222_us_71:
		next_state = LEGUP_F_main_BB_for_body222_us_72;
LEGUP_F_main_BB_for_body222_us_72:
		next_state = LEGUP_F_main_BB_for_body222_us_73;
LEGUP_F_main_BB_for_body222_us_73:
	if ((fsm_stall == 1'd0) && (main_for_body222_us_cmp224_us_reg == 1'd1))
		next_state = LEGUP_F_main_BB_if_then226_us_74;
	else if ((fsm_stall == 1'd0) && (main_for_body222_us_cmp224_us_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc291_us_78;
LEGUP_F_main_BB_for_body222_us_preheader_70:
		next_state = LEGUP_F_main_BB_for_body222_us_71;
LEGUP_F_main_BB_for_body300_84:
		next_state = LEGUP_F_main_BB_for_body300_85;
LEGUP_F_main_BB_for_body300_85:
		next_state = LEGUP_F_main_BB_for_body_i_86;
LEGUP_F_main_BB_for_body300_preheader_83:
		next_state = LEGUP_F_main_BB_for_body300_84;
LEGUP_F_main_BB_for_body6_i_90:
		next_state = LEGUP_F_main_BB_for_body_i_i_91;
LEGUP_F_main_BB_for_body_i_86:
		next_state = LEGUP_F_main_BB_for_body_i_87;
LEGUP_F_main_BB_for_body_i_87:
	if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond2_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_end_i_88;
	else if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond2_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_i_86;
LEGUP_F_main_BB_for_body_i_i_91:
		next_state = LEGUP_F_main_BB_for_body_i_i_92;
LEGUP_F_main_BB_for_body_i_i_92:
	if ((fsm_stall == 1'd0) && (main_for_body_i_i_cmp1_i_i == 1'd1))
		next_state = LEGUP_F_main_BB_land_lhs_true_i_i_93;
	else if ((fsm_stall == 1'd0) && (main_for_body_i_i_cmp1_i_i == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc_i_i_95;
LEGUP_F_main_BB_for_cond171_preheader_44:
		next_state = LEGUP_F_main_BB_for_cond171_preheader_45;
LEGUP_F_main_BB_for_cond171_preheader_45:
		next_state = LEGUP_F_main_BB_for_body173_46;
LEGUP_F_main_BB_for_cond186_preheader_53:
		next_state = LEGUP_F_main_BB_for_cond186_preheader_54;
LEGUP_F_main_BB_for_cond186_preheader_54:
		next_state = LEGUP_F_main_BB_for_body188_55;
LEGUP_F_main_BB_for_cond186_preheader_preheader_52:
		next_state = LEGUP_F_main_BB_for_cond186_preheader_53;
LEGUP_F_main_BB_for_cond220_preheader_68:
		next_state = LEGUP_F_main_BB_for_cond220_preheader_69;
LEGUP_F_main_BB_for_cond220_preheader_69:
	if ((fsm_stall == 1'd0) && (main_for_cond220_preheader_cmp223_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_body222_us_preheader_70;
	else if ((fsm_stall == 1'd0) && (main_for_cond220_preheader_cmp223_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc291_8_120;
LEGUP_F_main_BB_for_cond220_preheader_preheader_67:
		next_state = LEGUP_F_main_BB_for_cond220_preheader_68;
LEGUP_F_main_BB_for_end342_119:
		next_state = LEGUP_0;
LEGUP_F_main_BB_for_end342_loopexit1_118:
		next_state = LEGUP_F_main_BB_for_end342_119;
LEGUP_F_main_BB_for_end342_loopexit_117:
		next_state = LEGUP_F_main_BB_for_end342_119;
LEGUP_F_main_BB_for_end_i_88:
		next_state = LEGUP_F_main_BB_for_end_i_89;
LEGUP_F_main_BB_for_end_i_89:
		next_state = LEGUP_F_main_BB_for_body6_i_90;
LEGUP_F_main_BB_for_inc178_51:
	if ((fsm_stall == 1'd0) && (main_for_inc178_exitcond12 == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond186_preheader_preheader_52;
	else if ((fsm_stall == 1'd0) && (main_for_inc178_exitcond12 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond171_preheader_44;
LEGUP_F_main_BB_for_inc195_59:
	if ((fsm_stall == 1'd0) && (main_for_inc195_exitcond == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc198_60;
	else if ((fsm_stall == 1'd0) && (main_for_inc195_exitcond == 1'd0))
		next_state = LEGUP_F_main_BB_for_body188_55;
LEGUP_F_main_BB_for_inc198_60:
	if ((fsm_stall == 1'd0) && (main_for_inc198_exitcond10 == 1'd1))
		next_state = LEGUP_F_main_BB_for_body203_preheader_61;
	else if ((fsm_stall == 1'd0) && (main_for_inc198_exitcond10 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond186_preheader_53;
LEGUP_F_main_BB_for_inc214_66:
	if ((fsm_stall == 1'd0) && (main_for_inc214_exitcond9 == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond220_preheader_preheader_67;
	else if ((fsm_stall == 1'd0) && (main_for_inc214_exitcond9 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body203_62;
LEGUP_F_main_BB_for_inc28_i_106:
	if ((fsm_stall == 1'd0) && (main_for_inc28_i_exitcond4 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc31_i_107;
	else if ((fsm_stall == 1'd0) && (main_for_inc28_i_exitcond4 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body11_i_98;
LEGUP_F_main_BB_for_inc291_8_120:
		next_state = LEGUP_F_main_BB_for_inc291_8_121;
LEGUP_F_main_BB_for_inc291_8_121:
		next_state = LEGUP_F_main_BB_for_inc291_8_122;
LEGUP_F_main_BB_for_inc291_8_122:
		next_state = LEGUP_F_main_BB_for_inc291_8_123;
LEGUP_F_main_BB_for_inc291_8_123:
		next_state = LEGUP_F_main_BB_for_inc291_8_124;
LEGUP_F_main_BB_for_inc291_8_124:
		next_state = LEGUP_F_main_BB_for_inc291_8_125;
LEGUP_F_main_BB_for_inc291_8_125:
		next_state = LEGUP_F_main_BB_for_inc291_8_126;
LEGUP_F_main_BB_for_inc291_8_126:
		next_state = LEGUP_F_main_BB_for_inc291_8_127;
LEGUP_F_main_BB_for_inc291_8_127:
		next_state = LEGUP_F_main_BB_for_inc291_8_128;
LEGUP_F_main_BB_for_inc291_8_128:
		next_state = LEGUP_F_main_BB_for_inc291_8_129;
LEGUP_F_main_BB_for_inc291_8_129:
		next_state = LEGUP_F_main_BB_for_inc294_82;
LEGUP_F_main_BB_for_inc291_us_78:
		next_state = LEGUP_F_main_BB_for_inc291_us_79;
LEGUP_F_main_BB_for_inc291_us_79:
		next_state = LEGUP_F_main_BB_for_inc291_us_80;
LEGUP_F_main_BB_for_inc291_us_80:
	if ((fsm_stall == 1'd0) && (main_for_inc291_us_exitcond6_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc294_loopexit_81;
	else if ((fsm_stall == 1'd0) && (main_for_inc291_us_exitcond6_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body222_us_71;
LEGUP_F_main_BB_for_inc294_82:
	if ((fsm_stall == 1'd0) && (main_for_inc294_exitcond7 == 1'd1))
		next_state = LEGUP_F_main_BB_for_body300_preheader_83;
	else if ((fsm_stall == 1'd0) && (main_for_inc294_exitcond7 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond220_preheader_68;
LEGUP_F_main_BB_for_inc294_loopexit_81:
		next_state = LEGUP_F_main_BB_for_inc294_82;
LEGUP_F_main_BB_for_inc31_i_107:
	if ((fsm_stall == 1'd0) && (main_for_inc31_i_exitcond5 == 1'd1))
		next_state = LEGUP_F_main_BB_dijkstra_exit_108;
	else if ((fsm_stall == 1'd0) && (main_for_inc31_i_exitcond5 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body6_i_90;
LEGUP_F_main_BB_for_inc340_116:
	if ((fsm_stall == 1'd0) && (main_for_inc340_cmp298 == 1'd1))
		next_state = LEGUP_F_main_BB_for_body300_84;
	else if ((fsm_stall == 1'd0) && (main_for_inc340_cmp298 == 1'd0))
		next_state = LEGUP_F_main_BB_for_end342_loopexit1_118;
LEGUP_F_main_BB_for_inc340_loopexit_115:
		next_state = LEGUP_F_main_BB_for_inc340_116;
LEGUP_F_main_BB_for_inc_50:
	if ((fsm_stall == 1'd0) && (main_for_inc_exitcond11 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc178_51;
	else if ((fsm_stall == 1'd0) && (main_for_inc_exitcond11 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body173_46;
LEGUP_F_main_BB_for_inc_i_i_95:
	if ((fsm_stall == 1'd0) && (main_for_inc_i_i_exitcond3 == 1'd1))
		next_state = LEGUP_F_main_BB_minDistance_exit_i_96;
	else if ((fsm_stall == 1'd0) && (main_for_inc_i_i_exitcond3 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_i_i_91;
LEGUP_F_main_BB_if_end313_111:
		next_state = LEGUP_F_main_BB_if_end313_112;
LEGUP_F_main_BB_if_end313_112:
	if ((fsm_stall == 1'd0) && (main_if_end313_and320425 == 1'd1))
		next_state = LEGUP_F_main_BB_if_then322_113;
	else if ((fsm_stall == 1'd0) && (main_if_end313_and320425 == 1'd0))
		next_state = LEGUP_F_main_BB_for_end342_loopexit_117;
LEGUP_F_main_BB_if_end313_preheader_110:
		next_state = LEGUP_F_main_BB_if_end313_111;
LEGUP_F_main_BB_if_then192_57:
		next_state = LEGUP_F_main_BB_if_then192_58;
LEGUP_F_main_BB_if_then192_58:
		next_state = LEGUP_F_main_BB_for_inc195_59;
LEGUP_F_main_BB_if_then226_us_74:
		next_state = LEGUP_F_main_BB_if_then226_us_75;
LEGUP_F_main_BB_if_then226_us_75:
		next_state = LEGUP_F_main_BB_if_then226_us_76;
LEGUP_F_main_BB_if_then226_us_76:
		next_state = LEGUP_F_main_BB_if_then226_us_77;
LEGUP_F_main_BB_if_then226_us_77:
		next_state = LEGUP_F_main_BB_for_inc291_us_78;
LEGUP_F_main_BB_if_then322_113:
		next_state = LEGUP_F_main_BB_if_then322_114;
LEGUP_F_main_BB_if_then322_114:
	if ((fsm_stall == 1'd0) && (main_if_then322_cmp310 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc340_loopexit_115;
	else if ((fsm_stall == 1'd0) && (main_if_then322_cmp310 == 1'd0))
		next_state = LEGUP_F_main_BB_if_end313_111;
LEGUP_F_main_BB_if_then_48:
		next_state = LEGUP_F_main_BB_if_then_49;
LEGUP_F_main_BB_if_then_49:
		next_state = LEGUP_F_main_BB_for_inc_50;
LEGUP_F_main_BB_if_then_i_104:
		next_state = LEGUP_F_main_BB_if_then_i_105;
LEGUP_F_main_BB_if_then_i_105:
		next_state = LEGUP_F_main_BB_for_inc28_i_106;
LEGUP_F_main_BB_land_lhs_true16_i_102:
		next_state = LEGUP_F_main_BB_land_lhs_true16_i_103;
LEGUP_F_main_BB_land_lhs_true16_i_103:
	if ((fsm_stall == 1'd0) && (main_land_lhs_true16_i_cmp21_i == 1'd1))
		next_state = LEGUP_F_main_BB_if_then_i_104;
	else if ((fsm_stall == 1'd0) && (main_land_lhs_true16_i_cmp21_i == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc28_i_106;
LEGUP_F_main_BB_land_lhs_true_i_100:
		next_state = LEGUP_F_main_BB_land_lhs_true_i_101;
LEGUP_F_main_BB_land_lhs_true_i_101:
	if ((fsm_stall == 1'd0) && (main_land_lhs_true_i_tobool15_i == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc28_i_106;
	else if ((fsm_stall == 1'd0) && (main_land_lhs_true_i_tobool15_i == 1'd0))
		next_state = LEGUP_F_main_BB_land_lhs_true16_i_102;
LEGUP_F_main_BB_land_lhs_true_i_i_93:
		next_state = LEGUP_F_main_BB_land_lhs_true_i_i_94;
LEGUP_F_main_BB_land_lhs_true_i_i_94:
		next_state = LEGUP_F_main_BB_for_inc_i_i_95;
LEGUP_F_main_BB_minDistance_exit_i_96:
		next_state = LEGUP_F_main_BB_minDistance_exit_i_97;
LEGUP_F_main_BB_minDistance_exit_i_97:
		next_state = LEGUP_F_main_BB_for_body11_i_98;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
assign main_entry_vla1422_sub = 1'd0;
assign main_entry_vla421_sub = 1'd0;
assign main_entry_arrayidx3 = (1'd0 + (4 * 32'd1));
assign main_entry_arrayidx4 = (1'd0 + (4 * 32'd1));
assign main_entry_arrayidx5 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx5_reg <= main_entry_arrayidx5;
	end
end
assign main_entry_arrayidx6 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx6_reg <= main_entry_arrayidx6;
	end
end
assign main_entry_arrayidx7 = (1'd0 + (4 * 32'd3));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx7_reg <= main_entry_arrayidx7;
	end
end
assign main_entry_arrayidx8 = (1'd0 + (4 * 32'd3));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx8_reg <= main_entry_arrayidx8;
	end
end
assign main_entry_arrayidx9 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx9_reg <= main_entry_arrayidx9;
	end
end
assign main_entry_arrayidx10 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx10_reg <= main_entry_arrayidx10;
	end
end
assign main_entry_arrayidx11 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx11_reg <= main_entry_arrayidx11;
	end
end
assign main_entry_arrayidx12 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx12_reg <= main_entry_arrayidx12;
	end
end
assign main_entry_arrayidx13 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx13_reg <= main_entry_arrayidx13;
	end
end
assign main_entry_arrayidx14 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx14_reg <= main_entry_arrayidx14;
	end
end
assign main_entry_arrayidx15 = (1'd0 + (4 * 32'd7));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx15_reg <= main_entry_arrayidx15;
	end
end
assign main_entry_arrayidx16 = (1'd0 + (4 * 32'd7));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx16_reg <= main_entry_arrayidx16;
	end
end
assign main_entry_arrayidx17 = (1'd0 + (4 * 32'd8));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx17_reg <= main_entry_arrayidx17;
	end
end
assign main_entry_arrayidx18 = (1'd0 + (4 * 32'd8));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx18_reg <= main_entry_arrayidx18;
	end
end
assign main_entry_arrayidx19 = (1'd0 + (4 * 32'd9));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx19_reg <= main_entry_arrayidx19;
	end
end
assign main_entry_arrayidx20 = (1'd0 + (4 * 32'd9));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx20_reg <= main_entry_arrayidx20;
	end
end
assign main_entry_arrayidx21 = (1'd0 + (4 * 32'd10));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx21_reg <= main_entry_arrayidx21;
	end
end
assign main_entry_arrayidx22 = (1'd0 + (4 * 32'd10));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx22_reg <= main_entry_arrayidx22;
	end
end
assign main_entry_arrayidx23 = (1'd0 + (4 * 32'd11));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx23_reg <= main_entry_arrayidx23;
	end
end
assign main_entry_arrayidx24 = (1'd0 + (4 * 32'd11));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx24_reg <= main_entry_arrayidx24;
	end
end
assign main_entry_arrayidx25 = (1'd0 + (4 * 32'd12));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx25_reg <= main_entry_arrayidx25;
	end
end
assign main_entry_arrayidx26 = (1'd0 + (4 * 32'd12));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx26_reg <= main_entry_arrayidx26;
	end
end
assign main_entry_arrayidx27 = (1'd0 + (4 * 32'd13));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx27_reg <= main_entry_arrayidx27;
	end
end
assign main_entry_arrayidx28 = (1'd0 + (4 * 32'd13));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx28_reg <= main_entry_arrayidx28;
	end
end
assign main_entry_arrayidx29 = (1'd0 + (4 * 32'd14));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx29_reg <= main_entry_arrayidx29;
	end
end
assign main_entry_arrayidx30 = (1'd0 + (4 * 32'd14));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx30_reg <= main_entry_arrayidx30;
	end
end
assign main_entry_arrayidx31 = (1'd0 + (4 * 32'd15));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx31_reg <= main_entry_arrayidx31;
	end
end
assign main_entry_arrayidx32 = (1'd0 + (4 * 32'd15));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx32_reg <= main_entry_arrayidx32;
	end
end
assign main_entry_arrayidx33 = (1'd0 + (4 * 32'd16));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx33_reg <= main_entry_arrayidx33;
	end
end
assign main_entry_arrayidx34 = (1'd0 + (4 * 32'd16));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx34_reg <= main_entry_arrayidx34;
	end
end
assign main_entry_arrayidx35 = (1'd0 + (4 * 32'd17));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx35_reg <= main_entry_arrayidx35;
	end
end
assign main_entry_arrayidx36 = (1'd0 + (4 * 32'd17));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx36_reg <= main_entry_arrayidx36;
	end
end
assign main_entry_arrayidx37 = (1'd0 + (4 * 32'd18));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx37_reg <= main_entry_arrayidx37;
	end
end
assign main_entry_arrayidx38 = (1'd0 + (4 * 32'd18));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx38_reg <= main_entry_arrayidx38;
	end
end
assign main_entry_arrayidx39 = (1'd0 + (4 * 32'd19));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx39_reg <= main_entry_arrayidx39;
	end
end
assign main_entry_arrayidx40 = (1'd0 + (4 * 32'd19));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx40_reg <= main_entry_arrayidx40;
	end
end
assign main_entry_arrayidx41 = (1'd0 + (4 * 32'd20));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx41_reg <= main_entry_arrayidx41;
	end
end
assign main_entry_arrayidx42 = (1'd0 + (4 * 32'd20));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx42_reg <= main_entry_arrayidx42;
	end
end
assign main_entry_arrayidx43 = (1'd0 + (4 * 32'd21));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx43_reg <= main_entry_arrayidx43;
	end
end
assign main_entry_arrayidx44 = (1'd0 + (4 * 32'd21));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx44_reg <= main_entry_arrayidx44;
	end
end
assign main_entry_arrayidx45 = (1'd0 + (4 * 32'd22));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx45_reg <= main_entry_arrayidx45;
	end
end
assign main_entry_arrayidx46 = (1'd0 + (4 * 32'd22));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx46_reg <= main_entry_arrayidx46;
	end
end
assign main_entry_arrayidx47 = (1'd0 + (4 * 32'd23));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx47_reg <= main_entry_arrayidx47;
	end
end
assign main_entry_arrayidx48 = (1'd0 + (4 * 32'd23));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx48_reg <= main_entry_arrayidx48;
	end
end
assign main_entry_arrayidx49 = (1'd0 + (4 * 32'd24));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx49_reg <= main_entry_arrayidx49;
	end
end
assign main_entry_arrayidx50 = (1'd0 + (4 * 32'd24));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx50_reg <= main_entry_arrayidx50;
	end
end
assign main_entry_arrayidx51 = (1'd0 + (4 * 32'd25));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx51_reg <= main_entry_arrayidx51;
	end
end
assign main_entry_arrayidx52 = (1'd0 + (4 * 32'd25));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx52_reg <= main_entry_arrayidx52;
	end
end
assign main_entry_arrayidx53 = (1'd0 + (4 * 32'd26));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx53_reg <= main_entry_arrayidx53;
	end
end
assign main_entry_arrayidx54 = (1'd0 + (4 * 32'd26));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx54_reg <= main_entry_arrayidx54;
	end
end
assign main_entry_arrayidx55 = (1'd0 + (4 * 32'd27));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx55_reg <= main_entry_arrayidx55;
	end
end
assign main_entry_arrayidx56 = (1'd0 + (4 * 32'd27));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx56_reg <= main_entry_arrayidx56;
	end
end
assign main_entry_arrayidx57 = (1'd0 + (4 * 32'd28));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx57_reg <= main_entry_arrayidx57;
	end
end
assign main_entry_arrayidx58 = (1'd0 + (4 * 32'd28));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx58_reg <= main_entry_arrayidx58;
	end
end
assign main_entry_arrayidx59 = (1'd0 + (4 * 32'd29));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx59_reg <= main_entry_arrayidx59;
	end
end
assign main_entry_arrayidx60 = (1'd0 + (4 * 32'd29));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx60_reg <= main_entry_arrayidx60;
	end
end
assign main_entry_arrayidx61 = (1'd0 + (4 * 32'd30));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx61_reg <= main_entry_arrayidx61;
	end
end
assign main_entry_arrayidx62 = (1'd0 + (4 * 32'd30));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx62_reg <= main_entry_arrayidx62;
	end
end
assign main_entry_arrayidx63 = (1'd0 + (4 * 32'd31));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx63_reg <= main_entry_arrayidx63;
	end
end
assign main_entry_arrayidx64 = (1'd0 + (4 * 32'd31));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx64_reg <= main_entry_arrayidx64;
	end
end
assign main_entry_arrayidx65 = (1'd0 + (4 * 32'd32));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx65_reg <= main_entry_arrayidx65;
	end
end
assign main_entry_arrayidx66 = (1'd0 + (4 * 32'd32));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx66_reg <= main_entry_arrayidx66;
	end
end
assign main_entry_arrayidx67 = (1'd0 + (4 * 32'd33));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx67_reg <= main_entry_arrayidx67;
	end
end
assign main_entry_arrayidx68 = (1'd0 + (4 * 32'd33));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx68_reg <= main_entry_arrayidx68;
	end
end
assign main_entry_arrayidx69 = (1'd0 + (4 * 32'd34));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx69_reg <= main_entry_arrayidx69;
	end
end
assign main_entry_arrayidx70 = (1'd0 + (4 * 32'd34));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx70_reg <= main_entry_arrayidx70;
	end
end
assign main_entry_arrayidx71 = (1'd0 + (4 * 32'd35));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx71_reg <= main_entry_arrayidx71;
	end
end
assign main_entry_arrayidx72 = (1'd0 + (4 * 32'd35));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx72_reg <= main_entry_arrayidx72;
	end
end
assign main_entry_arrayidx73 = (1'd0 + (4 * 32'd36));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx73_reg <= main_entry_arrayidx73;
	end
end
assign main_entry_arrayidx74 = (1'd0 + (4 * 32'd36));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx74_reg <= main_entry_arrayidx74;
	end
end
assign main_entry_arrayidx75 = (1'd0 + (4 * 32'd37));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx75_reg <= main_entry_arrayidx75;
	end
end
assign main_entry_arrayidx76 = (1'd0 + (4 * 32'd37));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx76_reg <= main_entry_arrayidx76;
	end
end
assign main_entry_arrayidx77 = (1'd0 + (4 * 32'd38));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx77_reg <= main_entry_arrayidx77;
	end
end
assign main_entry_arrayidx78 = (1'd0 + (4 * 32'd38));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx78_reg <= main_entry_arrayidx78;
	end
end
assign main_entry_arrayidx79 = (1'd0 + (4 * 32'd39));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx79_reg <= main_entry_arrayidx79;
	end
end
assign main_entry_arrayidx80 = (1'd0 + (4 * 32'd39));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx80_reg <= main_entry_arrayidx80;
	end
end
assign main_entry_arrayidx81 = (1'd0 + (4 * 32'd40));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx81_reg <= main_entry_arrayidx81;
	end
end
assign main_entry_arrayidx82 = (1'd0 + (4 * 32'd40));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx82_reg <= main_entry_arrayidx82;
	end
end
assign main_entry_arrayidx83 = (1'd0 + (4 * 32'd41));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx83_reg <= main_entry_arrayidx83;
	end
end
assign main_entry_arrayidx84 = (1'd0 + (4 * 32'd41));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx84_reg <= main_entry_arrayidx84;
	end
end
assign main_entry_arrayidx85 = (1'd0 + (4 * 32'd42));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx85_reg <= main_entry_arrayidx85;
	end
end
assign main_entry_arrayidx86 = (1'd0 + (4 * 32'd42));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx86_reg <= main_entry_arrayidx86;
	end
end
assign main_entry_arrayidx87 = (1'd0 + (4 * 32'd43));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx87_reg <= main_entry_arrayidx87;
	end
end
assign main_entry_arrayidx88 = (1'd0 + (4 * 32'd43));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx88_reg <= main_entry_arrayidx88;
	end
end
assign main_entry_arrayidx89 = (1'd0 + (4 * 32'd44));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx89_reg <= main_entry_arrayidx89;
	end
end
assign main_entry_arrayidx90 = (1'd0 + (4 * 32'd44));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx90_reg <= main_entry_arrayidx90;
	end
end
assign main_entry_arrayidx91 = (1'd0 + (4 * 32'd45));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx91_reg <= main_entry_arrayidx91;
	end
end
assign main_entry_arrayidx92 = (1'd0 + (4 * 32'd45));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx92_reg <= main_entry_arrayidx92;
	end
end
assign main_entry_arrayidx93 = (1'd0 + (4 * 32'd46));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx93_reg <= main_entry_arrayidx93;
	end
end
assign main_entry_arrayidx94 = (1'd0 + (4 * 32'd46));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx94_reg <= main_entry_arrayidx94;
	end
end
assign main_entry_arrayidx95 = (1'd0 + (4 * 32'd47));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx95_reg <= main_entry_arrayidx95;
	end
end
assign main_entry_arrayidx96 = (1'd0 + (4 * 32'd47));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx96_reg <= main_entry_arrayidx96;
	end
end
assign main_entry_arrayidx97 = (1'd0 + (4 * 32'd48));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx97_reg <= main_entry_arrayidx97;
	end
end
assign main_entry_arrayidx98 = (1'd0 + (4 * 32'd48));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx98_reg <= main_entry_arrayidx98;
	end
end
assign main_entry_arrayidx99 = (1'd0 + (4 * 32'd49));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx99_reg <= main_entry_arrayidx99;
	end
end
assign main_entry_arrayidx100 = (1'd0 + (4 * 32'd49));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx100_reg <= main_entry_arrayidx100;
	end
end
assign main_entry_arrayidx101 = (1'd0 + (4 * 32'd50));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx101_reg <= main_entry_arrayidx101;
	end
end
assign main_entry_arrayidx102 = (1'd0 + (4 * 32'd50));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx102_reg <= main_entry_arrayidx102;
	end
end
assign main_entry_arrayidx103 = (1'd0 + (4 * 32'd51));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx103_reg <= main_entry_arrayidx103;
	end
end
assign main_entry_arrayidx104 = (1'd0 + (4 * 32'd51));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx104_reg <= main_entry_arrayidx104;
	end
end
assign main_entry_arrayidx105 = (1'd0 + (4 * 32'd52));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx105_reg <= main_entry_arrayidx105;
	end
end
assign main_entry_arrayidx106 = (1'd0 + (4 * 32'd52));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx106_reg <= main_entry_arrayidx106;
	end
end
assign main_entry_arrayidx107 = (1'd0 + (4 * 32'd53));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx107_reg <= main_entry_arrayidx107;
	end
end
assign main_entry_arrayidx108 = (1'd0 + (4 * 32'd53));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx108_reg <= main_entry_arrayidx108;
	end
end
assign main_entry_arrayidx109 = (1'd0 + (4 * 32'd54));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx109_reg <= main_entry_arrayidx109;
	end
end
assign main_entry_arrayidx110 = (1'd0 + (4 * 32'd54));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx110_reg <= main_entry_arrayidx110;
	end
end
assign main_entry_arrayidx111 = (1'd0 + (4 * 32'd55));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx111_reg <= main_entry_arrayidx111;
	end
end
assign main_entry_arrayidx112 = (1'd0 + (4 * 32'd55));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx112_reg <= main_entry_arrayidx112;
	end
end
assign main_entry_arrayidx113 = (1'd0 + (4 * 32'd56));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx113_reg <= main_entry_arrayidx113;
	end
end
assign main_entry_arrayidx114 = (1'd0 + (4 * 32'd56));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx114_reg <= main_entry_arrayidx114;
	end
end
assign main_entry_arrayidx115 = (1'd0 + (4 * 32'd57));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx115_reg <= main_entry_arrayidx115;
	end
end
assign main_entry_arrayidx116 = (1'd0 + (4 * 32'd57));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx116_reg <= main_entry_arrayidx116;
	end
end
assign main_entry_arrayidx117 = (1'd0 + (4 * 32'd58));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx117_reg <= main_entry_arrayidx117;
	end
end
assign main_entry_arrayidx118 = (1'd0 + (4 * 32'd58));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx118_reg <= main_entry_arrayidx118;
	end
end
assign main_entry_arrayidx119 = (1'd0 + (4 * 32'd59));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx119_reg <= main_entry_arrayidx119;
	end
end
assign main_entry_arrayidx120 = (1'd0 + (4 * 32'd59));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx120_reg <= main_entry_arrayidx120;
	end
end
assign main_entry_arrayidx121 = (1'd0 + (4 * 32'd60));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx121_reg <= main_entry_arrayidx121;
	end
end
assign main_entry_arrayidx122 = (1'd0 + (4 * 32'd60));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx122_reg <= main_entry_arrayidx122;
	end
end
assign main_entry_arrayidx123 = (1'd0 + (4 * 32'd61));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx123_reg <= main_entry_arrayidx123;
	end
end
assign main_entry_arrayidx124 = (1'd0 + (4 * 32'd61));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx124_reg <= main_entry_arrayidx124;
	end
end
assign main_entry_arrayidx125 = (1'd0 + (4 * 32'd62));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx125_reg <= main_entry_arrayidx125;
	end
end
assign main_entry_arrayidx126 = (1'd0 + (4 * 32'd62));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx126_reg <= main_entry_arrayidx126;
	end
end
assign main_entry_arrayidx127 = (1'd0 + (4 * 32'd63));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx127_reg <= main_entry_arrayidx127;
	end
end
assign main_entry_arrayidx128 = (1'd0 + (4 * 32'd63));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx128_reg <= main_entry_arrayidx128;
	end
end
assign main_entry_arrayidx129 = (1'd0 + (4 * 32'd64));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx129_reg <= main_entry_arrayidx129;
	end
end
assign main_entry_arrayidx130 = (1'd0 + (4 * 32'd64));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx130_reg <= main_entry_arrayidx130;
	end
end
assign main_entry_arrayidx131 = (1'd0 + (4 * 32'd65));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx131_reg <= main_entry_arrayidx131;
	end
end
assign main_entry_arrayidx132 = (1'd0 + (4 * 32'd65));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx132_reg <= main_entry_arrayidx132;
	end
end
assign main_entry_arrayidx133 = (1'd0 + (4 * 32'd66));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx133_reg <= main_entry_arrayidx133;
	end
end
assign main_entry_arrayidx134 = (1'd0 + (4 * 32'd66));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx134_reg <= main_entry_arrayidx134;
	end
end
assign main_entry_arrayidx135 = (1'd0 + (4 * 32'd67));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx135_reg <= main_entry_arrayidx135;
	end
end
assign main_entry_arrayidx136 = (1'd0 + (4 * 32'd67));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx136_reg <= main_entry_arrayidx136;
	end
end
assign main_entry_arrayidx137 = (1'd0 + (4 * 32'd68));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx137_reg <= main_entry_arrayidx137;
	end
end
assign main_entry_arrayidx138 = (1'd0 + (4 * 32'd68));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx138_reg <= main_entry_arrayidx138;
	end
end
assign main_entry_arrayidx139 = (1'd0 + (4 * 32'd69));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx139_reg <= main_entry_arrayidx139;
	end
end
assign main_entry_arrayidx140 = (1'd0 + (4 * 32'd69));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx140_reg <= main_entry_arrayidx140;
	end
end
assign main_entry_arrayidx141 = (1'd0 + (4 * 32'd70));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx141_reg <= main_entry_arrayidx141;
	end
end
assign main_entry_arrayidx142 = (1'd0 + (4 * 32'd70));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx142_reg <= main_entry_arrayidx142;
	end
end
assign main_entry_arrayidx143 = (1'd0 + (4 * 32'd71));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx143_reg <= main_entry_arrayidx143;
	end
end
assign main_entry_arrayidx144 = (1'd0 + (4 * 32'd71));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx144_reg <= main_entry_arrayidx144;
	end
end
assign main_entry_arrayidx145 = (1'd0 + (4 * 32'd72));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx145_reg <= main_entry_arrayidx145;
	end
end
assign main_entry_arrayidx146 = (1'd0 + (4 * 32'd72));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx146_reg <= main_entry_arrayidx146;
	end
end
assign main_entry_arrayidx147 = (1'd0 + (4 * 32'd73));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx147_reg <= main_entry_arrayidx147;
	end
end
assign main_entry_arrayidx148 = (1'd0 + (4 * 32'd73));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx148_reg <= main_entry_arrayidx148;
	end
end
assign main_entry_arrayidx149 = (1'd0 + (4 * 32'd74));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx149_reg <= main_entry_arrayidx149;
	end
end
assign main_entry_arrayidx150 = (1'd0 + (4 * 32'd74));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx150_reg <= main_entry_arrayidx150;
	end
end
assign main_entry_arrayidx151 = (1'd0 + (4 * 32'd75));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx151_reg <= main_entry_arrayidx151;
	end
end
assign main_entry_arrayidx152 = (1'd0 + (4 * 32'd75));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx152_reg <= main_entry_arrayidx152;
	end
end
assign main_entry_arrayidx153 = (1'd0 + (4 * 32'd76));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx153_reg <= main_entry_arrayidx153;
	end
end
assign main_entry_arrayidx154 = (1'd0 + (4 * 32'd76));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx154_reg <= main_entry_arrayidx154;
	end
end
assign main_entry_arrayidx155 = (1'd0 + (4 * 32'd77));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx155_reg <= main_entry_arrayidx155;
	end
end
assign main_entry_arrayidx156 = (1'd0 + (4 * 32'd77));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx156_reg <= main_entry_arrayidx156;
	end
end
assign main_entry_arrayidx157 = (1'd0 + (4 * 32'd78));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx157_reg <= main_entry_arrayidx157;
	end
end
assign main_entry_arrayidx158 = (1'd0 + (4 * 32'd78));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx158_reg <= main_entry_arrayidx158;
	end
end
assign main_entry_arrayidx159 = (1'd0 + (4 * 32'd79));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx159_reg <= main_entry_arrayidx159;
	end
end
assign main_entry_arrayidx160 = (1'd0 + (4 * 32'd79));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx160_reg <= main_entry_arrayidx160;
	end
end
assign main_entry_arrayidx161 = (1'd0 + (4 * 32'd80));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx161_reg <= main_entry_arrayidx161;
	end
end
assign main_entry_arrayidx162 = (1'd0 + (4 * 32'd80));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx162_reg <= main_entry_arrayidx162;
	end
end
assign main_entry_arrayidx163 = (1'd0 + (4 * 32'd81));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx163_reg <= main_entry_arrayidx163;
	end
end
assign main_entry_arrayidx164 = (1'd0 + (4 * 32'd81));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx164_reg <= main_entry_arrayidx164;
	end
end
assign main_entry_arrayidx165 = (1'd0 + (4 * 32'd82));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx165_reg <= main_entry_arrayidx165;
	end
end
assign main_entry_arrayidx166 = (1'd0 + (4 * 32'd82));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx166_reg <= main_entry_arrayidx166;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_entry_43) & (fsm_stall == 1'd0))) begin
		main_for_cond171_preheader_j169_0444 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc178_51) & (fsm_stall == 1'd0)) & (main_for_inc178_exitcond12 == 1'd0))) */ begin
		main_for_cond171_preheader_j169_0444 = main_for_inc178_4;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_entry_43) & (fsm_stall == 1'd0))) begin
		main_for_cond171_preheader_j169_0444_reg <= main_for_cond171_preheader_j169_0444;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc178_51) & (fsm_stall == 1'd0)) & (main_for_inc178_exitcond12 == 1'd0))) begin
		main_for_cond171_preheader_j169_0444_reg <= main_for_cond171_preheader_j169_0444;
	end
end
always @(*) begin
		main_for_cond171_preheader_arrayidx174 = (1'd0 + (4 * {25'd0,main_for_cond171_preheader_j169_0444_reg}));
end
always @(*) begin
		main_for_cond171_preheader_arrayidx177 = (1'd0 + (4 * {25'd0,main_for_cond171_preheader_j169_0444_reg}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond171_preheader_44)) begin
		main_for_cond171_preheader_arrayidx177_reg <= main_for_cond171_preheader_arrayidx177;
	end
end
always @(*) begin
		main_for_cond171_preheader_0 = main_entry_vla421_out_b;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond171_preheader_45)) begin
		main_for_cond171_preheader_0_reg <= main_for_cond171_preheader_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond171_preheader_45) & (fsm_stall == 1'd0))) begin
		main_for_body173_1 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_50) & (fsm_stall == 1'd0)) & (main_for_inc_exitcond11 == 1'd0))) */ begin
		main_for_body173_1 = main_for_inc_3;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond171_preheader_45) & (fsm_stall == 1'd0))) begin
		main_for_body173_1_reg <= main_for_body173_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_50) & (fsm_stall == 1'd0)) & (main_for_inc_exitcond11 == 1'd0))) begin
		main_for_body173_1_reg <= main_for_body173_1;
	end
end
always @(*) begin
		main_for_body173_arrayidx175 = (1'd0 + (4 * main_for_body173_1_reg));
end
always @(*) begin
		main_for_body173_2 = main_grid_out_a;
end
always @(*) begin
		main_for_body173_cmp176 = (main_for_cond171_preheader_0_reg == main_for_body173_2);
end
always @(*) begin
		main_for_inc_3 = (main_for_body173_1_reg + 32'd1);
end
always @(*) begin
		main_for_inc_exitcond11 = (main_for_inc_3 == 32'd81);
end
always @(*) begin
		main_for_inc178_4 = ({1'd0,main_for_cond171_preheader_j169_0444_reg} + 32'd1);
end
always @(*) begin
		main_for_inc178_exitcond12 = (main_for_inc178_4 == 32'd83);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond186_preheader_preheader_52) & (fsm_stall == 1'd0))) begin
		main_for_cond186_preheader_j181_0442 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc198_60) & (fsm_stall == 1'd0)) & (main_for_inc198_exitcond10 == 1'd0))) */ begin
		main_for_cond186_preheader_j181_0442 = main_for_inc198_9;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond186_preheader_preheader_52) & (fsm_stall == 1'd0))) begin
		main_for_cond186_preheader_j181_0442_reg <= main_for_cond186_preheader_j181_0442;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc198_60) & (fsm_stall == 1'd0)) & (main_for_inc198_exitcond10 == 1'd0))) begin
		main_for_cond186_preheader_j181_0442_reg <= main_for_cond186_preheader_j181_0442;
	end
end
always @(*) begin
		main_for_cond186_preheader_arrayidx189 = (1'd0 + (4 * {25'd0,main_for_cond186_preheader_j181_0442_reg}));
end
always @(*) begin
		main_for_cond186_preheader_arrayidx193 = (1'd0 + (4 * {25'd0,main_for_cond186_preheader_j181_0442_reg}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond186_preheader_53)) begin
		main_for_cond186_preheader_arrayidx193_reg <= main_for_cond186_preheader_arrayidx193;
	end
end
always @(*) begin
		main_for_cond186_preheader_5 = main_entry_vla1422_out_b;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond186_preheader_54)) begin
		main_for_cond186_preheader_5_reg <= main_for_cond186_preheader_5;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond186_preheader_54) & (fsm_stall == 1'd0))) begin
		main_for_body188_6 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc195_59) & (fsm_stall == 1'd0)) & (main_for_inc195_exitcond == 1'd0))) */ begin
		main_for_body188_6 = main_for_inc195_8;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond186_preheader_54) & (fsm_stall == 1'd0))) begin
		main_for_body188_6_reg <= main_for_body188_6;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc195_59) & (fsm_stall == 1'd0)) & (main_for_inc195_exitcond == 1'd0))) begin
		main_for_body188_6_reg <= main_for_body188_6;
	end
end
always @(*) begin
		main_for_body188_arrayidx190 = (1'd0 + (4 * main_for_body188_6_reg));
end
always @(*) begin
		main_for_body188_7 = main_grid_out_a;
end
always @(*) begin
		main_for_body188_cmp191 = (main_for_cond186_preheader_5_reg == main_for_body188_7);
end
always @(*) begin
		main_for_inc195_8 = (main_for_body188_6_reg + 32'd1);
end
always @(*) begin
		main_for_inc195_exitcond = (main_for_inc195_8 == 32'd81);
end
always @(*) begin
		main_for_inc198_9 = ({1'd0,main_for_cond186_preheader_j181_0442_reg} + 32'd1);
end
always @(*) begin
		main_for_inc198_exitcond10 = (main_for_inc198_9 == 32'd83);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body203_preheader_61) & (fsm_stall == 1'd0))) begin
		main_for_body203_i_0440 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc214_66) & (fsm_stall == 1'd0)) & (main_for_inc214_exitcond9 == 1'd0))) */ begin
		main_for_body203_i_0440 = main_for_inc214_11;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body203_preheader_61) & (fsm_stall == 1'd0))) begin
		main_for_body203_i_0440_reg <= main_for_body203_i_0440;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc214_66) & (fsm_stall == 1'd0)) & (main_for_inc214_exitcond9 == 1'd0))) begin
		main_for_body203_i_0440_reg <= main_for_body203_i_0440;
	end
end
always @(*) begin
		main_for_body203_arrayidx204 = (1'd0 + (4 * {25'd0,main_for_body203_i_0440_reg}));
end
always @(*) begin
		main_for_body203_arrayidx205 = (1'd0 + (4 * {25'd0,main_for_body203_i_0440_reg}));
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body203_63) & (fsm_stall == 1'd0))) begin
		main_for_body208_j_0439 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body208_65) & (fsm_stall == 1'd0)) & (main_for_body208_exitcond8_reg == 1'd0))) */ begin
		main_for_body208_j_0439 = main_for_body208_10_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body203_63) & (fsm_stall == 1'd0))) begin
		main_for_body208_j_0439_reg <= main_for_body208_j_0439;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body208_65) & (fsm_stall == 1'd0)) & (main_for_body208_exitcond8_reg == 1'd0))) begin
		main_for_body208_j_0439_reg <= main_for_body208_j_0439;
	end
end
always @(*) begin
		main_for_body208_arrayidx210 = (1'd0 + ((324 * {25'd0,main_for_body203_i_0440_reg}) + (4 * main_for_body208_j_0439_reg)));
end
always @(*) begin
		main_for_body208_10 = (main_for_body208_j_0439_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body208_64)) begin
		main_for_body208_10_reg <= main_for_body208_10;
	end
end
always @(*) begin
		main_for_body208_exitcond8 = (main_for_body208_10 == 32'd81);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body208_64)) begin
		main_for_body208_exitcond8_reg <= main_for_body208_exitcond8;
	end
end
always @(*) begin
		main_for_inc214_11 = ({1'd0,main_for_body203_i_0440_reg} + 32'd1);
end
always @(*) begin
		main_for_inc214_exitcond9 = (main_for_inc214_11 == 32'd81);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond220_preheader_preheader_67) & (fsm_stall == 1'd0))) begin
		main_for_cond220_preheader_12 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc294_82) & (fsm_stall == 1'd0)) & (main_for_inc294_exitcond7 == 1'd0))) */ begin
		main_for_cond220_preheader_12 = main_for_inc294_25;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond220_preheader_preheader_67) & (fsm_stall == 1'd0))) begin
		main_for_cond220_preheader_12_reg <= main_for_cond220_preheader_12;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc294_82) & (fsm_stall == 1'd0)) & (main_for_inc294_exitcond7 == 1'd0))) begin
		main_for_cond220_preheader_12_reg <= main_for_cond220_preheader_12;
	end
end
always @(*) begin
		main_for_cond220_preheader_bit_select13 = main_for_cond220_preheader_12_reg_width_extended[30:0];
end
always @(*) begin
		main_for_cond220_preheader_bit_select9 = main_for_cond220_preheader_12_reg_width_extended[23:0];
end
always @(*) begin
		main_for_cond220_preheader_bit_select7 = main_for_cond220_preheader_12_reg_width_extended[22:0];
end
always @(*) begin
		main_for_cond220_preheader_sr_negate = (32'd0 - {1'd0,main_for_cond220_preheader_12_reg});
end
always @(*) begin
		main_for_cond220_preheader_bit_select11 = main_for_cond220_preheader_sr_negate_width_extended[26:0];
end
always @(*) begin
		main_for_cond220_preheader_bit_concat14 = {main_for_cond220_preheader_bit_select13[30:0], main_for_cond220_preheader_bit_concat14_bit_select_operand_2};
end
always @(*) begin
		main_for_cond220_preheader_bit_concat12 = {main_for_cond220_preheader_bit_select11[26:0], main_for_cond220_preheader_bit_concat12_bit_select_operand_2[4:0]};
end
always @(*) begin
		main_for_cond220_preheader_bit_concat10 = {main_for_cond220_preheader_bit_select9[23:0], main_for_cond220_preheader_bit_concat10_bit_select_operand_2[7:0]};
end
always @(*) begin
		main_for_cond220_preheader_bit_concat8 = {main_for_cond220_preheader_bit_select7[22:0], main_for_cond220_preheader_bit_concat8_bit_select_operand_2[8:0]};
end
always @(*) begin
		main_for_cond220_preheader_sr_add = (main_for_cond220_preheader_bit_concat14 + main_for_cond220_preheader_bit_concat12);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_68)) begin
		main_for_cond220_preheader_sr_add_reg <= main_for_cond220_preheader_sr_add;
	end
end
always @(*) begin
		main_for_cond220_preheader_sr_add16 = (main_for_cond220_preheader_bit_concat10 + main_for_cond220_preheader_bit_concat8);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_68)) begin
		main_for_cond220_preheader_sr_add16_reg <= main_for_cond220_preheader_sr_add16;
	end
end
always @(*) begin
		main_for_cond220_preheader_sr_add17 = (main_for_cond220_preheader_sr_add_reg + main_for_cond220_preheader_sr_add16_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_69)) begin
		main_for_cond220_preheader_sr_add17_reg <= main_for_cond220_preheader_sr_add17;
	end
end
always @(*) begin
		main_for_cond220_preheader_bit_select5 = main_for_cond220_preheader_sr_add17[31:1];
end
always @(*) begin
		main_for_cond220_preheader_13 = (main_for_cond220_preheader_sr_add17 + 32'd9);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_69)) begin
		main_for_cond220_preheader_13_reg <= main_for_cond220_preheader_13;
	end
end
always @(*) begin
		main_for_cond220_preheader_bit_concat6 = {main_for_cond220_preheader_bit_select5[30:0], main_for_cond220_preheader_bit_concat6_bit_select_operand_2};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_69)) begin
		main_for_cond220_preheader_bit_concat6_reg <= main_for_cond220_preheader_bit_concat6;
	end
end
always @(*) begin
		main_for_cond220_preheader_14 = (main_for_cond220_preheader_sr_add17 + 32'd2);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_69)) begin
		main_for_cond220_preheader_14_reg <= main_for_cond220_preheader_14;
	end
end
always @(*) begin
		main_for_cond220_preheader_15 = (main_for_cond220_preheader_sr_add17 + 32'd3);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_69)) begin
		main_for_cond220_preheader_15_reg <= main_for_cond220_preheader_15;
	end
end
always @(*) begin
		main_for_cond220_preheader_16 = (main_for_cond220_preheader_sr_add17 + 32'd4);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_69)) begin
		main_for_cond220_preheader_16_reg <= main_for_cond220_preheader_16;
	end
end
always @(*) begin
		main_for_cond220_preheader_17 = (main_for_cond220_preheader_sr_add17 + 32'd5);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_69)) begin
		main_for_cond220_preheader_17_reg <= main_for_cond220_preheader_17;
	end
end
always @(*) begin
		main_for_cond220_preheader_18 = (main_for_cond220_preheader_sr_add17 + 32'd6);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_69)) begin
		main_for_cond220_preheader_18_reg <= main_for_cond220_preheader_18;
	end
end
always @(*) begin
		main_for_cond220_preheader_19 = (main_for_cond220_preheader_sr_add17 + 32'd7);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_69)) begin
		main_for_cond220_preheader_19_reg <= main_for_cond220_preheader_19;
	end
end
always @(*) begin
		main_for_cond220_preheader_cmp223 = ($signed({27'd0,main_for_cond220_preheader_cmp223_op0_temp}) < $signed({26'd0,main_for_cond220_preheader_cmp223_op1_temp}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond220_preheader_68)) begin
		main_for_cond220_preheader_cmp223_reg <= main_for_cond220_preheader_cmp223;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body222_us_preheader_70) & (fsm_stall == 1'd0))) begin
		main_for_body222_us_20 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc291_us_80) & (fsm_stall == 1'd0)) & (main_for_inc291_us_exitcond6_reg == 1'd0))) */ begin
		main_for_body222_us_20 = main_for_inc291_us_24_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body222_us_preheader_70) & (fsm_stall == 1'd0))) begin
		main_for_body222_us_20_reg <= main_for_body222_us_20;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc291_us_80) & (fsm_stall == 1'd0)) & (main_for_inc291_us_exitcond6_reg == 1'd0))) begin
		main_for_body222_us_20_reg <= main_for_body222_us_20;
	end
end
always @(*) begin
		main_for_body222_us_bit_select3 = main_for_body222_us_20_reg[30:0];
end
always @(*) begin
		main_for_body222_us_bit_select1 = main_for_body222_us_20_reg[27:0];
end
always @(*) begin
		main_for_body222_us_bit_select = main_for_body222_us_20_reg[25:0];
end
always @(*) begin
		main_for_body222_us_bit_concat4 = {main_for_body222_us_bit_select3[30:0], main_for_body222_us_bit_concat4_bit_select_operand_2};
end
always @(*) begin
		main_for_body222_us_bit_concat2 = {main_for_body222_us_bit_select1[27:0], main_for_body222_us_bit_concat2_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body222_us_bit_concat = {main_for_body222_us_bit_select[25:0], main_for_body222_us_bit_concat_bit_select_operand_2[5:0]};
end
always @(*) begin
		main_for_body222_us_sr_add21 = (main_for_body222_us_bit_concat4 + main_for_body222_us_bit_concat2);
end
always @(*) begin
		main_for_body222_us_sr_add22 = (main_for_body222_us_bit_concat + main_for_body222_us_sr_add21);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body222_us_71)) begin
		main_for_body222_us_sr_add22_reg <= main_for_body222_us_sr_add22;
	end
end
always @(*) begin
		main_for_body222_us_21 = (main_for_cond220_preheader_13_reg + main_for_body222_us_sr_add22_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body222_us_72)) begin
		main_for_body222_us_21_reg <= main_for_body222_us_21;
	end
end
always @(*) begin
		main_for_body222_us_arrayidx262_us = (1'd0 + (4 * main_for_body222_us_21_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body222_us_73)) begin
		main_for_body222_us_arrayidx262_us_reg <= main_for_body222_us_arrayidx262_us;
	end
end
always @(*) begin
		main_for_body222_us_22 = (main_for_cond220_preheader_sr_add17_reg + main_for_body222_us_sr_add22_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body222_us_72)) begin
		main_for_body222_us_22_reg <= main_for_body222_us_22;
	end
end
always @(*) begin
		main_for_body222_us_arrayidx269_us = (1'd0 + ((324 * 32'd9) + (4 * main_for_body222_us_22_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body222_us_73)) begin
		main_for_body222_us_arrayidx269_us_reg <= main_for_body222_us_arrayidx269_us;
	end
end
always @(*) begin
		main_for_body222_us_cmp224_us = ($signed(main_for_body222_us_20_reg) < $signed({26'd0,main_for_body222_us_cmp224_us_op1_temp}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body222_us_71)) begin
		main_for_body222_us_cmp224_us_reg <= main_for_body222_us_cmp224_us;
	end
end
always @(*) begin
		main_if_then226_us_23 = (main_for_cond220_preheader_bit_concat6_reg + main_for_body222_us_sr_add22_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_then226_us_74)) begin
		main_if_then226_us_23_reg <= main_if_then226_us_23;
	end
end
always @(*) begin
		main_if_then226_us_arrayidx231_us = (1'd0 + (4 * main_if_then226_us_23_reg));
end
always @(*) begin
		main_if_then226_us_arrayidx238_us = (1'd0 + ((324 * 32'd1) + (4 * main_for_body222_us_22_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_then226_us_74)) begin
		main_if_then226_us_arrayidx238_us_reg <= main_if_then226_us_arrayidx238_us;
	end
end
always @(*) begin
		main_for_inc291_us_24 = (main_for_body222_us_20_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_us_78)) begin
		main_for_inc291_us_24_reg <= main_for_inc291_us_24;
	end
end
always @(*) begin
		main_for_inc291_us_exitcond6 = (main_for_inc291_us_24 == 32'd9);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_us_78)) begin
		main_for_inc291_us_exitcond6_reg <= main_for_inc291_us_exitcond6;
	end
end
always @(*) begin
		main_for_inc294_25 = ({1'd0,main_for_cond220_preheader_12_reg} + 32'd1);
end
always @(*) begin
		main_for_inc294_exitcond7 = (main_for_inc294_25 == 32'd9);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body300_preheader_83) & (fsm_stall == 1'd0))) begin
		main_for_body300_i_2435 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc340_116) & (fsm_stall == 1'd0)) & (main_for_inc340_cmp298 == 1'd1))) */ begin
		main_for_body300_i_2435 = main_for_body300_inc341_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body300_preheader_83) & (fsm_stall == 1'd0))) begin
		main_for_body300_i_2435_reg <= main_for_body300_i_2435;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc340_116) & (fsm_stall == 1'd0)) & (main_for_inc340_cmp298 == 1'd1))) begin
		main_for_body300_i_2435_reg <= main_for_body300_i_2435;
	end
end
always @(*) begin
		main_for_body300_arrayidx301 = (1'd0 + (4 * {25'd0,main_for_body300_i_2435_reg}));
end
always @(*) begin
		main_for_body300_arrayidx302 = (1'd0 + (4 * {25'd0,main_for_body300_i_2435_reg}));
end
always @(*) begin
		main_for_body300_inc341 = ({1'd0,main_for_body300_i_2435_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body300_84)) begin
		main_for_body300_inc341_reg <= main_for_body300_inc341;
	end
end
always @(*) begin
		main_for_body300_26 = main_entry_vla167423_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body300_85)) begin
		main_for_body300_26_reg <= main_for_body300_26;
	end
end
always @(*) begin
		main_for_body300_27 = main_entry_vla168424_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body300_85)) begin
		main_for_body300_27_reg <= main_for_body300_27;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body300_85) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_057_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body_i_87) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond2_reg == 1'd0))) */ begin
		main_for_body_i_i_057_i = main_for_body_i_28_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body300_85) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_057_i_reg <= main_for_body_i_i_057_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_87) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond2_reg == 1'd0))) begin
		main_for_body_i_i_057_i_reg <= main_for_body_i_i_057_i;
	end
end
always @(*) begin
		main_for_body_i_arrayidx1_i = (1'd0 + (4 * main_for_body_i_i_057_i_reg));
end
always @(*) begin
		main_for_body_i_arrayidx2_i = (1'd0 + (4 * main_for_body_i_i_057_i_reg));
end
always @(*) begin
		main_for_body_i_28 = (main_for_body_i_i_057_i_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_86)) begin
		main_for_body_i_28_reg <= main_for_body_i_28;
	end
end
always @(*) begin
		main_for_body_i_exitcond2 = (main_for_body_i_28 == 32'd81);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_86)) begin
		main_for_body_i_exitcond2_reg <= main_for_body_i_exitcond2;
	end
end
always @(*) begin
		main_for_end_i_arrayidx_i = (1'd0 + (4 * main_for_body300_26_reg));
end
always @(*) begin
		main_for_end_i_arrayidx3_i = (1'd0 + (4 * main_for_body300_26_reg));
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_end_i_89) & (fsm_stall == 1'd0))) begin
		main_for_body6_i_count_056_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc31_i_107) & (fsm_stall == 1'd0)) & (main_for_inc31_i_exitcond5 == 1'd0))) */ begin
		main_for_body6_i_count_056_i = main_for_inc31_i_38;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_end_i_89) & (fsm_stall == 1'd0))) begin
		main_for_body6_i_count_056_i_reg <= main_for_body6_i_count_056_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc31_i_107) & (fsm_stall == 1'd0)) & (main_for_inc31_i_exitcond5 == 1'd0))) begin
		main_for_body6_i_count_056_i_reg <= main_for_body6_i_count_056_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_90) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_29 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_95) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond3 == 1'd0))) */ begin
		main_for_body_i_i_29 = main_for_inc_i_i_32;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_90) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_29_reg <= main_for_body_i_i_29;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_95) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond3 == 1'd0))) begin
		main_for_body_i_i_29_reg <= main_for_body_i_i_29;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_90) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_index_012_i_i = 0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_95) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond3 == 1'd0))) */ begin
		main_for_body_i_i_min_index_012_i_i = main_for_inc_i_i_min_index_1_i_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_90) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_index_012_i_i_reg <= main_for_body_i_i_min_index_012_i_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_95) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond3 == 1'd0))) begin
		main_for_body_i_i_min_index_012_i_i_reg <= main_for_body_i_i_min_index_012_i_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_90) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_011_i_i = 32'd2147483647;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_95) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond3 == 1'd0))) */ begin
		main_for_body_i_i_min_011_i_i = main_for_inc_i_i_min_1_i_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_90) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_011_i_i_reg <= main_for_body_i_i_min_011_i_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_95) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond3 == 1'd0))) begin
		main_for_body_i_i_min_011_i_i_reg <= main_for_body_i_i_min_011_i_i;
	end
end
always @(*) begin
		main_for_body_i_i_arrayidx_i_i = (1'd0 + (4 * main_for_body_i_i_29_reg));
end
always @(*) begin
		main_for_body_i_i_30 = main_entry_sptSet_i_out_a;
end
always @(*) begin
		main_for_body_i_i_cmp1_i_i = (main_for_body_i_i_30 == 32'd0);
end
always @(*) begin
		main_land_lhs_true_i_i_arrayidx2_i_i = (1'd0 + (4 * main_for_body_i_i_29_reg));
end
always @(*) begin
		main_land_lhs_true_i_i_31 = main_entry_dist_i_out_a;
end
always @(*) begin
		main_land_lhs_true_i_i_cmp3_i_i = ($signed(main_land_lhs_true_i_i_31) > $signed(main_for_body_i_i_min_011_i_i_reg));
end
always @(*) begin
		main_land_lhs_true_i_i_min_0_i_i = (main_land_lhs_true_i_i_cmp3_i_i ? main_for_body_i_i_min_011_i_i_reg : main_land_lhs_true_i_i_31);
end
always @(*) begin
		main_land_lhs_true_i_i_min_index_0_v_0_i_i = (main_land_lhs_true_i_i_cmp3_i_i ? main_for_body_i_i_min_index_012_i_i_reg : main_for_body_i_i_29_reg);
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_92) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_1_i_i = main_for_body_i_i_min_011_i_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_94) & (fsm_stall == 1'd0))) */ begin
		main_for_inc_i_i_min_1_i_i = main_land_lhs_true_i_i_min_0_i_i;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_92) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_1_i_i_reg <= main_for_inc_i_i_min_1_i_i;
	end
	if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_94) & (fsm_stall == 1'd0))) begin
		main_for_inc_i_i_min_1_i_i_reg <= main_for_inc_i_i_min_1_i_i;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_92) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_index_1_i_i = main_for_body_i_i_min_index_012_i_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_94) & (fsm_stall == 1'd0))) */ begin
		main_for_inc_i_i_min_index_1_i_i = main_land_lhs_true_i_i_min_index_0_v_0_i_i;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_92) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_index_1_i_i_reg <= main_for_inc_i_i_min_index_1_i_i;
	end
	if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_94) & (fsm_stall == 1'd0))) begin
		main_for_inc_i_i_min_index_1_i_i_reg <= main_for_inc_i_i_min_index_1_i_i;
	end
end
always @(*) begin
		main_for_inc_i_i_32 = (main_for_body_i_i_29_reg + 32'd1);
end
always @(*) begin
		main_for_inc_i_i_exitcond3 = (main_for_inc_i_i_32 == 32'd81);
end
always @(*) begin
		main_minDistance_exit_i_arrayidx8_i = (1'd0 + (4 * main_for_inc_i_i_min_index_1_i_i_reg));
end
always @(*) begin
		main_minDistance_exit_i_arrayidx17_i = (1'd0 + (4 * main_for_inc_i_i_min_index_1_i_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_96)) begin
		main_minDistance_exit_i_arrayidx17_i_reg <= main_minDistance_exit_i_arrayidx17_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_minDistance_exit_i_97) & (fsm_stall == 1'd0))) begin
		main_for_body11_i_v_055_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc28_i_106) & (fsm_stall == 1'd0)) & (main_for_inc28_i_exitcond4 == 1'd0))) */ begin
		main_for_body11_i_v_055_i = main_for_inc28_i_37;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_minDistance_exit_i_97) & (fsm_stall == 1'd0))) begin
		main_for_body11_i_v_055_i_reg <= main_for_body11_i_v_055_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc28_i_106) & (fsm_stall == 1'd0)) & (main_for_inc28_i_exitcond4 == 1'd0))) begin
		main_for_body11_i_v_055_i_reg <= main_for_body11_i_v_055_i;
	end
end
always @(*) begin
		main_for_body11_i_arrayidx12_i = (1'd0 + (4 * main_for_body11_i_v_055_i_reg));
end
always @(*) begin
		main_for_body11_i_arrayidx20_i = (1'd0 + (4 * main_for_body11_i_v_055_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body11_i_98)) begin
		main_for_body11_i_arrayidx20_i_reg <= main_for_body11_i_arrayidx20_i;
	end
end
always @(*) begin
		main_for_body11_i_arrayidx22_i = (1'd0 + (4 * main_for_body11_i_v_055_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body11_i_98)) begin
		main_for_body11_i_arrayidx22_i_reg <= main_for_body11_i_arrayidx22_i;
	end
end
always @(*) begin
		main_for_body11_i_33 = main_entry_sptSet_i_out_a;
end
always @(*) begin
		main_for_body11_i_tobool_i = (main_for_body11_i_33 == 32'd0);
end
always @(*) begin
		main_land_lhs_true_i_arrayidx14_i = (1'd0 + ((324 * main_for_inc_i_i_min_index_1_i_i_reg) + (4 * main_for_body11_i_v_055_i_reg)));
end
always @(*) begin
		main_land_lhs_true_i_34 = main_entry_m_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_101)) begin
		main_land_lhs_true_i_34_reg <= main_land_lhs_true_i_34;
	end
end
always @(*) begin
		main_land_lhs_true_i_tobool15_i = (main_land_lhs_true_i_34 == 32'd0);
end
always @(*) begin
		main_land_lhs_true16_i_35 = main_entry_dist_i_out_a;
end
always @(*) begin
		main_land_lhs_true16_i_add_i = (main_land_lhs_true16_i_35 + main_land_lhs_true_i_34_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true16_i_103)) begin
		main_land_lhs_true16_i_add_i_reg <= main_land_lhs_true16_i_add_i;
	end
end
always @(*) begin
		main_land_lhs_true16_i_36 = main_entry_dist_i_out_b;
end
always @(*) begin
		main_land_lhs_true16_i_cmp21_i = ($signed(main_land_lhs_true16_i_add_i) < $signed(main_land_lhs_true16_i_36));
end
always @(*) begin
		main_for_inc28_i_37 = (main_for_body11_i_v_055_i_reg + 32'd1);
end
always @(*) begin
		main_for_inc28_i_exitcond4 = (main_for_inc28_i_37 == 32'd81);
end
always @(*) begin
		main_for_inc31_i_38 = (main_for_body6_i_count_056_i_reg + 32'd1);
end
always @(*) begin
		main_for_inc31_i_exitcond5 = (main_for_inc31_i_38 == 32'd80);
end
always @(*) begin
		main_dijkstra_exit_arrayidx309431 = (1'd0 + (4 * main_for_body300_27_reg));
end
always @(*) begin
		main_dijkstra_exit_39 = main_entry_parent_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_dijkstra_exit_109)) begin
		main_dijkstra_exit_39_reg <= main_dijkstra_exit_39;
	end
end
always @(*) begin
		main_dijkstra_exit_cmp310432 = (main_dijkstra_exit_39 == $signed(-32'd1));
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_end313_preheader_110) & (fsm_stall == 1'd0))) begin
		main_if_end313_40 = main_dijkstra_exit_39_reg;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_if_then322_114) & (fsm_stall == 1'd0)) & (main_if_then322_cmp310 == 1'd0))) */ begin
		main_if_end313_40 = main_if_then322_43;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_end313_preheader_110) & (fsm_stall == 1'd0))) begin
		main_if_end313_40_reg <= main_if_end313_40;
	end
	if ((((cur_state == LEGUP_F_main_BB_if_then322_114) & (fsm_stall == 1'd0)) & (main_if_then322_cmp310 == 1'd0))) begin
		main_if_end313_40_reg <= main_if_end313_40;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_end313_preheader_110) & (fsm_stall == 1'd0))) begin
		main_if_end313_origem_1434 = main_for_body300_27_reg;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_if_then322_114) & (fsm_stall == 1'd0)) & (main_if_then322_cmp310 == 1'd0))) */ begin
		main_if_end313_origem_1434 = main_if_end313_40_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_end313_preheader_110) & (fsm_stall == 1'd0))) begin
		main_if_end313_origem_1434_reg <= main_if_end313_origem_1434;
	end
	if ((((cur_state == LEGUP_F_main_BB_if_then322_114) & (fsm_stall == 1'd0)) & (main_if_then322_cmp310 == 1'd0))) begin
		main_if_end313_origem_1434_reg <= main_if_end313_origem_1434;
	end
end
always @(*) begin
		main_if_end313_arrayidx314 = (1'd0 + (4 * main_if_end313_40_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end313_111)) begin
		main_if_end313_arrayidx314_reg <= main_if_end313_arrayidx314;
	end
end
always @(*) begin
		main_if_end313_41 = main_entry_indice_s_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end313_112)) begin
		main_if_end313_41_reg <= main_if_end313_41;
	end
end
always @(*) begin
		main_if_end313_cmp315 = ($signed(main_if_end313_41) < $signed({27'd0,main_if_end313_cmp315_op1_temp}));
end
always @(*) begin
		main_if_end313_arrayidx317 = (1'd0 + (4 * main_if_end313_origem_1434_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end313_111)) begin
		main_if_end313_arrayidx317_reg <= main_if_end313_arrayidx317;
	end
end
always @(*) begin
		main_if_end313_42 = main_entry_indice_e_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end313_112)) begin
		main_if_end313_42_reg <= main_if_end313_42;
	end
end
always @(*) begin
		main_if_end313_cmp318 = ($signed(main_if_end313_42) < $signed({27'd0,main_if_end313_cmp318_op1_temp}));
end
always @(*) begin
		main_if_end313_and320425 = (main_if_end313_cmp315 & main_if_end313_cmp318);
end
always @(*) begin
		main_if_then322_add330 = (main_if_end313_42_reg + 32'd1);
end
always @(*) begin
		main_if_then322_add332 = (main_if_end313_41_reg + 32'd1);
end
always @(*) begin
		main_if_then322_arrayidx309 = (1'd0 + (4 * main_if_end313_40_reg));
end
always @(*) begin
		main_if_then322_43 = main_entry_parent_out_a;
end
always @(*) begin
		main_if_then322_cmp310 = (main_if_then322_43 == $signed(-32'd1));
end
always @(*) begin
		main_for_inc340_cmp298 = ($signed({23'd0,main_for_inc340_cmp298_op0_temp}) < $signed({23'd0,main_for_inc340_cmp298_op1_temp}));
end
always @(*) begin
		main_for_inc291_8_arrayidx287_1 = (1'd0 + ((324 * 32'd2) + (4 * main_for_cond220_preheader_bit_concat6_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx287_1_reg <= main_for_inc291_8_arrayidx287_1;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx280 = (1'd0 + (4 * main_for_cond220_preheader_bit_concat6_reg));
end
always @(*) begin
		main_for_inc291_8_arrayidx287 = (1'd0 + ((324 * 32'd1) + (4 * main_for_cond220_preheader_sr_add17_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx287_reg <= main_for_inc291_8_arrayidx287;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx287_7 = (1'd0 + ((324 * 32'd8) + (4 * main_for_cond220_preheader_19_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx287_7_reg <= main_for_inc291_8_arrayidx287_7;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx280_6 = (1'd0 + ((324 * 32'd6) + (4 * main_for_cond220_preheader_19_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx280_6_reg <= main_for_inc291_8_arrayidx280_6;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx287_6 = (1'd0 + ((324 * 32'd7) + (4 * main_for_cond220_preheader_18_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx287_6_reg <= main_for_inc291_8_arrayidx287_6;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx280_5 = (1'd0 + ((324 * 32'd5) + (4 * main_for_cond220_preheader_18_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx280_5_reg <= main_for_inc291_8_arrayidx280_5;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx287_5 = (1'd0 + ((324 * 32'd6) + (4 * main_for_cond220_preheader_17_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx287_5_reg <= main_for_inc291_8_arrayidx287_5;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx280_4 = (1'd0 + ((324 * 32'd4) + (4 * main_for_cond220_preheader_17_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx280_4_reg <= main_for_inc291_8_arrayidx280_4;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx287_4 = (1'd0 + ((324 * 32'd5) + (4 * main_for_cond220_preheader_16_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx287_4_reg <= main_for_inc291_8_arrayidx287_4;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx280_3 = (1'd0 + ((324 * 32'd3) + (4 * main_for_cond220_preheader_16_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx280_3_reg <= main_for_inc291_8_arrayidx280_3;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx287_3 = (1'd0 + ((324 * 32'd4) + (4 * main_for_cond220_preheader_15_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx287_3_reg <= main_for_inc291_8_arrayidx287_3;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx280_2 = (1'd0 + ((324 * 32'd2) + (4 * main_for_cond220_preheader_15_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx280_2_reg <= main_for_inc291_8_arrayidx280_2;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx287_2 = (1'd0 + ((324 * 32'd3) + (4 * main_for_cond220_preheader_14_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx287_2_reg <= main_for_inc291_8_arrayidx287_2;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx280_1 = (1'd0 + ((324 * 32'd1) + (4 * main_for_cond220_preheader_14_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_arrayidx280_1_reg <= main_for_inc291_8_arrayidx280_1;
	end
end
always @(*) begin
		main_for_inc291_8_44 = (main_for_cond220_preheader_sr_add17_reg + 32'd8);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_for_inc291_8_44_reg <= main_for_inc291_8_44;
	end
end
always @(*) begin
		main_for_inc291_8_arrayidx280_7 = (1'd0 + ((324 * 32'd7) + (4 * main_for_inc291_8_44_reg)));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_121)) begin
		main_for_inc291_8_arrayidx280_7_reg <= main_for_inc291_8_arrayidx280_7;
	end
end
always @(*) begin
	main_grid_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body173_46)) begin
		main_grid_address_a = (main_for_body173_arrayidx175 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body188_55)) begin
		main_grid_address_a = (main_for_body188_arrayidx190 >>> 3'd2);
	end
end
assign main_grid_address_b = 'dx;
always @(*) begin
	main_entry_dist_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_86)) begin
		main_entry_dist_i_address_a = (main_for_body_i_arrayidx1_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_end_i_88)) begin
		main_entry_dist_i_address_a = (main_for_end_i_arrayidx3_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_93)) begin
		main_entry_dist_i_address_a = (main_land_lhs_true_i_i_arrayidx2_i_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true16_i_102)) begin
		main_entry_dist_i_address_a = (main_minDistance_exit_i_arrayidx17_i_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_dist_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_86)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end_i_88)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_dist_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_86)) begin
		main_entry_dist_i_in_a = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end_i_88)) begin
		main_entry_dist_i_in_a = 32'd0;
	end
end
always @(*) begin
	main_entry_dist_i_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true16_i_102)) begin
		main_entry_dist_i_address_b = (main_for_body11_i_arrayidx20_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_104)) begin
		main_entry_dist_i_address_b = (main_for_body11_i_arrayidx20_i_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_dist_i_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_if_then_i_104)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_dist_i_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then_i_104)) begin
		main_entry_dist_i_in_b = main_land_lhs_true16_i_add_i_reg;
	end
end
always @(*) begin
	main_entry_sptSet_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_86)) begin
		main_entry_sptSet_i_address_a = (main_for_body_i_arrayidx2_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_i_91)) begin
		main_entry_sptSet_i_address_a = (main_for_body_i_i_arrayidx_i_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_96)) begin
		main_entry_sptSet_i_address_a = (main_minDistance_exit_i_arrayidx8_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body11_i_98)) begin
		main_entry_sptSet_i_address_a = (main_for_body11_i_arrayidx12_i >>> 3'd2);
	end
end
always @(*) begin
	main_entry_sptSet_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_86)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_96)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_sptSet_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_86)) begin
		main_entry_sptSet_i_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_96)) begin
		main_entry_sptSet_i_in_a = 32'd1;
	end
end
always @(*) begin
	main_entry_parent_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_end_i_88)) begin
		main_entry_parent_address_a = (main_for_end_i_arrayidx_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_104)) begin
		main_entry_parent_address_a = (main_for_body11_i_arrayidx22_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_dijkstra_exit_108)) begin
		main_entry_parent_address_a = (main_dijkstra_exit_arrayidx309431 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then322_113)) begin
		main_entry_parent_address_a = (main_if_then322_arrayidx309 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_parent_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_end_i_88)) begin
		main_entry_parent_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_104)) begin
		main_entry_parent_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_parent_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_end_i_88)) begin
		main_entry_parent_in_a = -32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_104)) begin
		main_entry_parent_in_a = main_for_inc_i_i_min_index_1_i_i_reg;
	end
end
always @(*) begin
	main_entry_m_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body208_64)) begin
		main_entry_m_address_a = (main_for_body208_arrayidx210 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then226_us_75)) begin
		main_entry_m_address_a = (main_if_then226_us_arrayidx231_us >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then226_us_76)) begin
		main_entry_m_address_a = (main_if_then226_us_arrayidx238_us_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_us_78)) begin
		main_entry_m_address_a = (main_for_body222_us_arrayidx262_us_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_us_79)) begin
		main_entry_m_address_a = (main_for_body222_us_arrayidx269_us_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_100)) begin
		main_entry_m_address_a = (main_land_lhs_true_i_arrayidx14_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_121)) begin
		main_entry_m_address_a = (main_for_inc291_8_arrayidx287_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_123)) begin
		main_entry_m_address_a = (main_for_inc291_8_arrayidx280_2_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_124)) begin
		main_entry_m_address_a = (main_for_inc291_8_arrayidx280_3_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_125)) begin
		main_entry_m_address_a = (main_for_inc291_8_arrayidx280_4_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_126)) begin
		main_entry_m_address_a = (main_for_inc291_8_arrayidx280_5_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_127)) begin
		main_entry_m_address_a = (main_for_inc291_8_arrayidx280_6_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_128)) begin
		main_entry_m_address_a = (main_for_inc291_8_arrayidx280_7_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_m_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body208_64)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then226_us_75)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then226_us_76)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_us_78)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_us_79)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_121)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_123)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_124)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_125)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_126)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_127)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_128)) begin
		main_entry_m_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_m_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body208_64)) begin
		main_entry_m_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then226_us_75)) begin
		main_entry_m_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then226_us_76)) begin
		main_entry_m_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_us_78)) begin
		main_entry_m_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_us_79)) begin
		main_entry_m_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_121)) begin
		main_entry_m_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_123)) begin
		main_entry_m_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_124)) begin
		main_entry_m_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_125)) begin
		main_entry_m_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_126)) begin
		main_entry_m_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_127)) begin
		main_entry_m_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_128)) begin
		main_entry_m_in_a = 32'd1;
	end
end
always @(*) begin
	main_entry_m_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_entry_m_address_b = (main_for_inc291_8_arrayidx280 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_121)) begin
		main_entry_m_address_b = (main_for_inc291_8_arrayidx280_1_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_122)) begin
		main_entry_m_address_b = (main_for_inc291_8_arrayidx287_1_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_123)) begin
		main_entry_m_address_b = (main_for_inc291_8_arrayidx287_2_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_124)) begin
		main_entry_m_address_b = (main_for_inc291_8_arrayidx287_3_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_125)) begin
		main_entry_m_address_b = (main_for_inc291_8_arrayidx287_4_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_126)) begin
		main_entry_m_address_b = (main_for_inc291_8_arrayidx287_5_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_127)) begin
		main_entry_m_address_b = (main_for_inc291_8_arrayidx287_6_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_128)) begin
		main_entry_m_address_b = (main_for_inc291_8_arrayidx287_7_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_m_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_entry_m_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_121)) begin
		main_entry_m_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_122)) begin
		main_entry_m_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_123)) begin
		main_entry_m_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_124)) begin
		main_entry_m_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_125)) begin
		main_entry_m_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_126)) begin
		main_entry_m_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_127)) begin
		main_entry_m_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_128)) begin
		main_entry_m_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_m_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_120)) begin
		main_entry_m_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_121)) begin
		main_entry_m_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_122)) begin
		main_entry_m_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_123)) begin
		main_entry_m_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_124)) begin
		main_entry_m_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_125)) begin
		main_entry_m_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_126)) begin
		main_entry_m_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_127)) begin
		main_entry_m_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc291_8_128)) begin
		main_entry_m_in_b = 32'd1;
	end
end
always @(*) begin
	main_entry_indice_e_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body203_62)) begin
		main_entry_indice_e_address_a = (main_for_body203_arrayidx204 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end313_111)) begin
		main_entry_indice_e_address_a = (main_if_end313_arrayidx317 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then322_113)) begin
		main_entry_indice_e_address_a = (main_if_end313_arrayidx317_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_indice_e_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body203_62)) begin
		main_entry_indice_e_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then322_113)) begin
		main_entry_indice_e_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_indice_e_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body203_62)) begin
		main_entry_indice_e_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then322_113)) begin
		main_entry_indice_e_in_a = main_if_then322_add330;
	end
end
always @(*) begin
	main_entry_indice_s_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body203_62)) begin
		main_entry_indice_s_address_a = (main_for_body203_arrayidx205 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end313_111)) begin
		main_entry_indice_s_address_a = (main_if_end313_arrayidx314 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then322_113)) begin
		main_entry_indice_s_address_a = (main_if_end313_arrayidx314_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_indice_s_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body203_62)) begin
		main_entry_indice_s_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then322_113)) begin
		main_entry_indice_s_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_indice_s_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body203_62)) begin
		main_entry_indice_s_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then322_113)) begin
		main_entry_indice_s_in_a = main_if_then322_add332;
	end
end
always @(*) begin
	main_entry_vla421_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla421_address_a = (main_entry_vla421_sub >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx5_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx9_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx13_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx17_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx21_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx25_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx29_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx33_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx37_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx41_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx45_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx49_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx53_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx57_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx61_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx65_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx69_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx73_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx77_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx81_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx85_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx89_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx93_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx97_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx101_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx105_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx109_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx113_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx117_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx121_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx125_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx129_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx133_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx137_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx141_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx145_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx149_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx153_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx157_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx161_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_42)) begin
		main_entry_vla421_address_a = (main_entry_arrayidx165_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla421_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_42)) begin
		main_entry_vla421_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla421_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla421_in_a = 32'd67;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla421_in_a = 32'd66;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla421_in_a = 32'd63;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla421_in_a = 32'd56;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla421_in_a = 32'd47;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla421_in_a = 32'd31;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla421_in_a = 32'd20;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla421_in_a = 32'd13;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla421_in_a = 32'd64;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla421_in_a = 32'd58;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla421_in_a = 32'd49;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla421_in_a = 32'd34;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla421_in_a = 32'd14;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla421_in_a = 32'd61;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla421_in_a = 32'd59;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla421_in_a = 32'd51;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla421_in_a = 32'd38;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla421_in_a = 32'd29;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla421_in_a = 32'd18;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla421_in_a = 32'd57;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla421_in_a = 32'd53;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla421_in_a = 32'd50;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla421_in_a = 32'd46;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla421_in_a = 32'd30;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla421_in_a = 32'd23;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla421_in_a = 32'd43;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla421_in_a = 32'd36;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla421_in_a = 32'd15;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla421_in_a = 32'd35;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla421_in_a = 32'd32;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla421_in_a = 32'd9;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla421_in_a = 32'd26;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla421_in_a = 32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla421_in_a = 32'd48;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla421_in_a = 32'd44;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla421_in_a = 32'd33;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla421_in_a = 32'd12;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla421_in_a = 32'd37;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla421_in_a = 32'd28;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla421_in_a = 32'd10;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla421_in_a = 32'd16;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_42)) begin
		main_entry_vla421_in_a = 32'd7;
	end
end
always @(*) begin
	main_entry_vla421_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx3 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx7_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx11_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx15_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx19_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx23_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx27_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx31_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx35_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx39_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx43_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx47_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx51_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx55_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx59_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx63_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx67_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx71_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx75_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx79_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx83_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx87_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx91_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx95_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx99_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx103_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx107_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx111_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx115_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx119_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx123_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx127_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx131_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx135_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx139_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx143_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx147_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx151_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx155_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx159_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla421_address_b = (main_entry_arrayidx163_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond171_preheader_44)) begin
		main_entry_vla421_address_b = (main_for_cond171_preheader_arrayidx174 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla421_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla421_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_vla421_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla421_in_b = 32'd66;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla421_in_b = 32'd65;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla421_in_b = 32'd60;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla421_in_b = 32'd52;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla421_in_b = 32'd40;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla421_in_b = 32'd20;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla421_in_b = 32'd8;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla421_in_b = 32'd64;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla421_in_b = 32'd62;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla421_in_b = 32'd54;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla421_in_b = 32'd42;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla421_in_b = 32'd25;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla421_in_b = 32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla421_in_b = 32'd61;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla421_in_b = 32'd55;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla421_in_b = 32'd45;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla421_in_b = 32'd29;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla421_in_b = 32'd19;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla421_in_b = 32'd6;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla421_in_b = 32'd57;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla421_in_b = 32'd53;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla421_in_b = 32'd50;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla421_in_b = 32'd39;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla421_in_b = 32'd30;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla421_in_b = 32'd11;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla421_in_b = 32'd43;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla421_in_b = 32'd27;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla421_in_b = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla421_in_b = 32'd35;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla421_in_b = 32'd21;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla421_in_b = 32'd26;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla421_in_b = 32'd17;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla421_in_b = 32'd48;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla421_in_b = 32'd44;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla421_in_b = 32'd41;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla421_in_b = 32'd24;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla421_in_b = 32'd37;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla421_in_b = 32'd28;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla421_in_b = 32'd22;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla421_in_b = 32'd16;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla421_in_b = 32'd7;
	end
end
always @(*) begin
	main_entry_vla1422_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1422_address_a = (main_entry_vla1422_sub >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx6_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx10_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx14_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx18_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx22_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx26_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx30_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx34_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx38_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx42_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx46_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx50_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx54_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx58_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx62_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx66_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx70_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx74_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx78_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx82_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx86_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx90_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx94_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx98_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx102_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx106_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx110_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx114_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx118_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx122_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx126_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx130_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx134_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx138_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx142_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx146_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx150_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx154_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx158_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx162_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_42)) begin
		main_entry_vla1422_address_a = (main_entry_arrayidx166_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla1422_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_42)) begin
		main_entry_vla1422_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla1422_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1422_in_a = 32'd66;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1422_in_a = 32'd65;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1422_in_a = 32'd60;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1422_in_a = 32'd52;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1422_in_a = 32'd40;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1422_in_a = 32'd20;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1422_in_a = 32'd8;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1422_in_a = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1422_in_a = 32'd62;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1422_in_a = 32'd54;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1422_in_a = 32'd42;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1422_in_a = 32'd25;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1422_in_a = 32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1422_in_a = 32'd57;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1422_in_a = 32'd55;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1422_in_a = 32'd45;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla1422_in_a = 32'd29;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla1422_in_a = 32'd19;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla1422_in_a = 32'd6;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla1422_in_a = 32'd53;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla1422_in_a = 32'd48;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla1422_in_a = 32'd46;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla1422_in_a = 32'd39;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla1422_in_a = 32'd19;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla1422_in_a = 32'd11;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla1422_in_a = 32'd35;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla1422_in_a = 32'd27;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla1422_in_a = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla1422_in_a = 32'd32;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla1422_in_a = 32'd21;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla1422_in_a = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla1422_in_a = 32'd15;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla1422_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla1422_in_a = 32'd42;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla1422_in_a = 32'd41;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla1422_in_a = 32'd24;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla1422_in_a = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla1422_in_a = 32'd27;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla1422_in_a = 32'd22;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla1422_in_a = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla1422_in_a = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_42)) begin
		main_entry_vla1422_in_a = 32'd1;
	end
end
always @(*) begin
	main_entry_vla1422_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx4 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx8_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx12_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx16_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx20_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx24_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx28_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx32_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx36_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx40_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx44_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx48_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx52_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx56_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx60_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx64_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx68_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx72_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx76_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx80_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx84_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx88_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx92_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx96_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx100_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx104_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx108_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx112_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx116_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx120_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx124_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx128_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx132_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx136_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx140_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx144_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx148_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx152_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx156_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx160_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla1422_address_b = (main_entry_arrayidx164_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond186_preheader_53)) begin
		main_entry_vla1422_address_b = (main_for_cond186_preheader_arrayidx189 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla1422_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla1422_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_vla1422_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1422_in_b = 32'd64;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1422_in_b = 32'd63;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1422_in_b = 32'd56;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1422_in_b = 32'd47;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1422_in_b = 32'd31;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1422_in_b = 32'd13;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1422_in_b = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1422_in_b = 32'd61;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1422_in_b = 32'd58;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1422_in_b = 32'd49;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1422_in_b = 32'd34;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1422_in_b = 32'd14;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1422_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1422_in_b = 32'd59;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1422_in_b = 32'd51;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1422_in_b = 32'd38;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_17)) begin
		main_entry_vla1422_in_b = 32'd18;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_18)) begin
		main_entry_vla1422_in_b = 32'd8;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_19)) begin
		main_entry_vla1422_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_20)) begin
		main_entry_vla1422_in_b = 32'd54;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_21)) begin
		main_entry_vla1422_in_b = 32'd50;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_22)) begin
		main_entry_vla1422_in_b = 32'd43;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_23)) begin
		main_entry_vla1422_in_b = 32'd30;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_24)) begin
		main_entry_vla1422_in_b = 32'd23;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_25)) begin
		main_entry_vla1422_in_b = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_26)) begin
		main_entry_vla1422_in_b = 32'd36;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_27)) begin
		main_entry_vla1422_in_b = 32'd15;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_28)) begin
		main_entry_vla1422_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_29)) begin
		main_entry_vla1422_in_b = 32'd26;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_30)) begin
		main_entry_vla1422_in_b = 32'd9;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_31)) begin
		main_entry_vla1422_in_b = 32'd17;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_32)) begin
		main_entry_vla1422_in_b = 32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_33)) begin
		main_entry_vla1422_in_b = 32'd44;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_34)) begin
		main_entry_vla1422_in_b = 32'd37;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_35)) begin
		main_entry_vla1422_in_b = 32'd33;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_36)) begin
		main_entry_vla1422_in_b = 32'd12;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_37)) begin
		main_entry_vla1422_in_b = 32'd28;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_38)) begin
		main_entry_vla1422_in_b = 32'd16;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_39)) begin
		main_entry_vla1422_in_b = 32'd10;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_40)) begin
		main_entry_vla1422_in_b = 32'd7;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_41)) begin
		main_entry_vla1422_in_b = 32'd2;
	end
end
always @(*) begin
	main_entry_vla167423_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then_48)) begin
		main_entry_vla167423_address_a = (main_for_cond171_preheader_arrayidx177_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body300_84)) begin
		main_entry_vla167423_address_a = (main_for_body300_arrayidx301 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla167423_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_if_then_48)) begin
		main_entry_vla167423_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla167423_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then_48)) begin
		main_entry_vla167423_in_a = main_for_body173_1_reg;
	end
end
always @(*) begin
	main_entry_vla168424_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then192_57)) begin
		main_entry_vla168424_address_a = (main_for_cond186_preheader_arrayidx193_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body300_84)) begin
		main_entry_vla168424_address_a = (main_for_body300_arrayidx302 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla168424_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_if_then192_57)) begin
		main_entry_vla168424_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla168424_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then192_57)) begin
		main_entry_vla168424_in_a = main_for_body188_6_reg;
	end
end
always @(*) begin
	main_for_cond220_preheader_12_reg_width_extended = {27'd0,main_for_cond220_preheader_12_reg};
end
always @(*) begin
	main_for_cond220_preheader_sr_negate_width_extended = {{22{main_for_cond220_preheader_sr_negate[4]}},main_for_cond220_preheader_sr_negate};
end
assign main_for_cond220_preheader_bit_concat14_bit_select_operand_2 = 1'd0;
assign main_for_cond220_preheader_bit_concat12_bit_select_operand_2 = 5'd0;
assign main_for_cond220_preheader_bit_concat10_bit_select_operand_2 = 8'd0;
assign main_for_cond220_preheader_bit_concat8_bit_select_operand_2 = 9'd0;
always @(*) begin
	main_for_cond220_preheader_cmp223_op0_temp = {1'd0,main_for_cond220_preheader_12_reg};
end
assign main_for_cond220_preheader_cmp223_op1_temp = 32'd8;
assign main_for_cond220_preheader_bit_concat6_bit_select_operand_2 = 1'd1;
assign main_for_body222_us_bit_concat4_bit_select_operand_2 = 1'd0;
assign main_for_body222_us_bit_concat2_bit_select_operand_2 = 4'd0;
assign main_for_body222_us_bit_concat_bit_select_operand_2 = 6'd0;
assign main_for_body222_us_cmp224_us_op1_temp = 32'd8;
assign main_if_end313_cmp315_op1_temp = 32'd4;
assign main_if_end313_cmp318_op1_temp = 32'd4;
always @(*) begin
	main_for_inc340_cmp298_op0_temp = {1'd0,main_for_body300_inc341_reg};
end
assign main_for_inc340_cmp298_op1_temp = 32'd83;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end342_119)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end342_119)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "Arria10",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module ram_single_port_intel
(
	clk,
	clken,
	address_a,
	wren_a,
	data_a,
	byteena_a,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
    .wren_a (wren_a),
    .data_a (data_a),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.operation_mode = "SINGLE_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "Arria10",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module rom_dual_port
(
	clk,
	clken,
	address_a,
	q_a,
	address_b,
	q_b
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  init_file = {`MEM_INIT_DIR, "UNUSED.mif"};
parameter  latency = 1;

input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
reg [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
reg [(width_b-1):0] q_b_wire;

(* ram_init_file = init_file *) reg [width_a-1:0] ram [numwords_a-1:0];

integer i;
/* synthesis translate_off */
ALTERA_MF_MEMORY_INITIALIZATION mem ();
reg [8*256:1] ram_ver_file;
initial begin
	if (init_file == {`MEM_INIT_DIR, "UNUSED.mif"})
    begin
		for (i = 0; i < numwords_a; i = i + 1)
			ram[i] = 0;
    end
	else
    begin
        // modelsim can't read .mif files directly. So use Altera function to
        // convert them to .ver files
        mem.convert_to_ver_file(init_file, width_a, ram_ver_file);
        $readmemh(ram_ver_file, ram);
    end
end
/* synthesis translate_on */

localparam input_latency = ((latency - 1) >> 1);
localparam output_latency = (latency - 1) - input_latency;
integer j;

reg [(widthad_a-1):0] address_a_reg[input_latency:0];
reg [(widthad_b-1):0] address_b_reg[input_latency:0];

always @(*)
begin
  address_a_reg[0] = address_a;
  address_b_reg[0] = address_b;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < input_latency; j=j+1)
   begin
       address_a_reg[j+1] <= address_a_reg[j];
       address_b_reg[j+1] <= address_b_reg[j];
   end
end

always @ (posedge clk)
if (clken)
begin
    q_a_wire <= ram[address_a_reg[input_latency]];
end

always @ (posedge clk)
if (clken)
begin
    q_b_wire <= ram[address_b_reg[input_latency]];
end


reg [(width_a-1):0] q_a_reg[output_latency:0];

always @(*)
begin
   q_a_reg[0] <= q_a_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_a_reg[j+1] <= q_a_reg[j];
   end
end

assign q_a = q_a_reg[output_latency];
reg [(width_b-1):0] q_b_reg[output_latency:0];

always @(*)
begin
   q_b_reg[0] <= q_b_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_b_reg[j+1] <= q_b_reg[j];
   end
end

assign q_b = q_b_reg[output_latency];

endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
