// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Fri May  8 21:46:26 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [6:0] LEGUP_0 = 7'd0;
parameter [6:0] LEGUP_F_main_BB_entry_1 = 7'd1;
parameter [6:0] LEGUP_F_main_BB_entry_2 = 7'd2;
parameter [6:0] LEGUP_F_main_BB_entry_3 = 7'd3;
parameter [6:0] LEGUP_F_main_BB_entry_4 = 7'd4;
parameter [6:0] LEGUP_F_main_BB_entry_5 = 7'd5;
parameter [6:0] LEGUP_F_main_BB_entry_6 = 7'd6;
parameter [6:0] LEGUP_F_main_BB_entry_7 = 7'd7;
parameter [6:0] LEGUP_F_main_BB_entry_8 = 7'd8;
parameter [6:0] LEGUP_F_main_BB_entry_9 = 7'd9;
parameter [6:0] LEGUP_F_main_BB_entry_10 = 7'd10;
parameter [6:0] LEGUP_F_main_BB_entry_11 = 7'd11;
parameter [6:0] LEGUP_F_main_BB_entry_12 = 7'd12;
parameter [6:0] LEGUP_F_main_BB_entry_13 = 7'd13;
parameter [6:0] LEGUP_F_main_BB_entry_14 = 7'd14;
parameter [6:0] LEGUP_F_main_BB_entry_15 = 7'd15;
parameter [6:0] LEGUP_F_main_BB_entry_16 = 7'd16;
parameter [6:0] LEGUP_F_main_BB_entry_17 = 7'd17;
parameter [6:0] LEGUP_F_main_BB_for_cond69_preheader_18 = 7'd18;
parameter [6:0] LEGUP_F_main_BB_for_cond69_preheader_19 = 7'd19;
parameter [6:0] LEGUP_F_main_BB_for_body71_20 = 7'd20;
parameter [6:0] LEGUP_F_main_BB_for_body71_21 = 7'd21;
parameter [6:0] LEGUP_F_main_BB_if_then_22 = 7'd22;
parameter [6:0] LEGUP_F_main_BB_if_then_23 = 7'd23;
parameter [6:0] LEGUP_F_main_BB_for_inc_24 = 7'd24;
parameter [6:0] LEGUP_F_main_BB_for_inc76_25 = 7'd25;
parameter [6:0] LEGUP_F_main_BB_for_cond84_preheader_preheader_26 = 7'd26;
parameter [6:0] LEGUP_F_main_BB_for_cond84_preheader_27 = 7'd27;
parameter [6:0] LEGUP_F_main_BB_for_cond84_preheader_28 = 7'd28;
parameter [6:0] LEGUP_F_main_BB_for_body86_29 = 7'd29;
parameter [6:0] LEGUP_F_main_BB_for_body86_30 = 7'd30;
parameter [6:0] LEGUP_F_main_BB_if_then90_31 = 7'd31;
parameter [6:0] LEGUP_F_main_BB_if_then90_32 = 7'd32;
parameter [6:0] LEGUP_F_main_BB_for_inc93_33 = 7'd33;
parameter [6:0] LEGUP_F_main_BB_for_inc96_34 = 7'd34;
parameter [6:0] LEGUP_F_main_BB_for_body101_preheader_35 = 7'd35;
parameter [6:0] LEGUP_F_main_BB_for_body101_36 = 7'd36;
parameter [6:0] LEGUP_F_main_BB_for_body101_37 = 7'd37;
parameter [6:0] LEGUP_F_main_BB_for_body106_38 = 7'd38;
parameter [6:0] LEGUP_F_main_BB_for_body106_39 = 7'd39;
parameter [6:0] LEGUP_F_main_BB_for_body106_40 = 7'd40;
parameter [6:0] LEGUP_F_main_BB_for_inc112_41 = 7'd41;
parameter [6:0] LEGUP_F_main_BB_for_cond118_preheader_preheader_42 = 7'd42;
parameter [6:0] LEGUP_F_main_BB_for_cond118_preheader_43 = 7'd43;
parameter [6:0] LEGUP_F_main_BB_for_cond118_preheader_44 = 7'd44;
parameter [6:0] LEGUP_F_main_BB_for_cond118_preheader_45 = 7'd45;
parameter [6:0] LEGUP_F_main_BB_for_cond118_preheader_46 = 7'd46;
parameter [6:0] LEGUP_F_main_BB_for_cond118_preheader_47 = 7'd47;
parameter [6:0] LEGUP_F_main_BB_for_inc192_48 = 7'd48;
parameter [6:0] LEGUP_F_main_BB_for_body198_preheader_49 = 7'd49;
parameter [6:0] LEGUP_F_main_BB_for_body198_50 = 7'd50;
parameter [6:0] LEGUP_F_main_BB_for_body198_51 = 7'd51;
parameter [6:0] LEGUP_F_main_BB_for_body_i_52 = 7'd52;
parameter [6:0] LEGUP_F_main_BB_for_body_i_53 = 7'd53;
parameter [6:0] LEGUP_F_main_BB_for_end_i_54 = 7'd54;
parameter [6:0] LEGUP_F_main_BB_for_end_i_55 = 7'd55;
parameter [6:0] LEGUP_F_main_BB_for_body6_i_56 = 7'd56;
parameter [6:0] LEGUP_F_main_BB_for_body_i_i_57 = 7'd57;
parameter [6:0] LEGUP_F_main_BB_for_body_i_i_58 = 7'd58;
parameter [6:0] LEGUP_F_main_BB_land_lhs_true_i_i_59 = 7'd59;
parameter [6:0] LEGUP_F_main_BB_land_lhs_true_i_i_60 = 7'd60;
parameter [6:0] LEGUP_F_main_BB_for_inc_i_i_61 = 7'd61;
parameter [6:0] LEGUP_F_main_BB_minDistance_exit_i_62 = 7'd62;
parameter [6:0] LEGUP_F_main_BB_minDistance_exit_i_63 = 7'd63;
parameter [6:0] LEGUP_F_main_BB_for_body11_i_64 = 7'd64;
parameter [6:0] LEGUP_F_main_BB_for_body11_i_65 = 7'd65;
parameter [6:0] LEGUP_F_main_BB_land_lhs_true_i_66 = 7'd66;
parameter [6:0] LEGUP_F_main_BB_land_lhs_true_i_67 = 7'd67;
parameter [6:0] LEGUP_F_main_BB_land_lhs_true_i_68 = 7'd68;
parameter [6:0] LEGUP_F_main_BB_land_lhs_true16_i_69 = 7'd69;
parameter [6:0] LEGUP_F_main_BB_land_lhs_true16_i_70 = 7'd70;
parameter [6:0] LEGUP_F_main_BB_if_then_i_71 = 7'd71;
parameter [6:0] LEGUP_F_main_BB_if_then_i_72 = 7'd72;
parameter [6:0] LEGUP_F_main_BB_for_inc28_i_73 = 7'd73;
parameter [6:0] LEGUP_F_main_BB_for_inc31_i_74 = 7'd74;
parameter [6:0] LEGUP_F_main_BB_dijkstra_exit_75 = 7'd75;
parameter [6:0] LEGUP_F_main_BB_dijkstra_exit_76 = 7'd76;
parameter [6:0] LEGUP_F_main_BB_if_end211_preheader_77 = 7'd77;
parameter [6:0] LEGUP_F_main_BB_if_end211_78 = 7'd78;
parameter [6:0] LEGUP_F_main_BB_if_end211_79 = 7'd79;
parameter [6:0] LEGUP_F_main_BB_if_then220_80 = 7'd80;
parameter [6:0] LEGUP_F_main_BB_if_then220_81 = 7'd81;
parameter [6:0] LEGUP_F_main_BB_for_inc238_loopexit_82 = 7'd82;
parameter [6:0] LEGUP_F_main_BB_for_inc238_83 = 7'd83;
parameter [6:0] LEGUP_F_main_BB_for_end240_loopexit_84 = 7'd84;
parameter [6:0] LEGUP_F_main_BB_for_end240_loopexit1_85 = 7'd85;
parameter [6:0] LEGUP_F_main_BB_for_end240_86 = 7'd86;
parameter [6:0] LEGUP_F_main_BB_for_inc189_5_87 = 7'd87;
parameter [6:0] LEGUP_F_main_BB_for_inc189_5_88 = 7'd88;
parameter [6:0] LEGUP_F_main_BB_for_inc189_5_89 = 7'd89;
parameter [6:0] LEGUP_F_main_BB_for_inc189_5_90 = 7'd90;
parameter [6:0] LEGUP_F_main_BB_for_inc189_5_91 = 7'd91;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_92 = 7'd92;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_93 = 7'd93;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_94 = 7'd94;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_95 = 7'd95;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_96 = 7'd96;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_97 = 7'd97;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_98 = 7'd98;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_99 = 7'd99;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_100 = 7'd100;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_101 = 7'd101;
parameter [6:0] LEGUP_F_main_BB_for_inc189_us_5_102 = 7'd102;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [6:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [6:0] next_state;
wire  fsm_stall;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_vla1320_sub;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_vla319_sub;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx3;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx4;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx5_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx6_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx7;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx7_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx8;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx8_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx9;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx9_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx10;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx10_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx11;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx11_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx12;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx12_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx13;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx13_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx14;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx14_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx15;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx15_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx16;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx16_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx17;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx17_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx18;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx18_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx19;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx19_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx20;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx20_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx21;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx21_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx22;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx22_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx23;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx23_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx24;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx24_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx25;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx25_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx26;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx26_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx27;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx27_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx28;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx28_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx29;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx29_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx30;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx30_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx31;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx31_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx32;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx32_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx33;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx33_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx34;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx34_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx35;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx35_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx36;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx36_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx37;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx37_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx38;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx38_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx39;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx39_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx40;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx40_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx41;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx41_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx42;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx42_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx43;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx43_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx44;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx44_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx45;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx45_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx46;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx46_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx47;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx47_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx48;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx48_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx49;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx49_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx50;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx50_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx51;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx51_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx52;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx52_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx53;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx53_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx54;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx54_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx55;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx55_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx56;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx56_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx57;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx57_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx58;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx58_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx59;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx59_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx60;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx60_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx61;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx61_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx62;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx62_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx63;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx63_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx64;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_arrayidx64_reg;
reg [5:0] main_for_cond69_preheader_j67_0342;
reg [5:0] main_for_cond69_preheader_j67_0342_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond69_preheader_arrayidx72;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond69_preheader_arrayidx75;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond69_preheader_arrayidx75_reg;
reg [31:0] main_for_cond69_preheader_0;
reg [31:0] main_for_cond69_preheader_0_reg;
reg [31:0] main_for_body71_1;
reg [31:0] main_for_body71_1_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body71_arrayidx73;
reg [31:0] main_for_body71_2;
reg  main_for_body71_cmp74;
reg [31:0] main_for_inc_3;
reg  main_for_inc_exitcond72;
reg [6:0] main_for_inc76_4;
reg  main_for_inc76_exitcond74;
reg [5:0] main_for_cond84_preheader_j79_0340;
reg [5:0] main_for_cond84_preheader_j79_0340_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond84_preheader_arrayidx87;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond84_preheader_arrayidx91;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond84_preheader_arrayidx91_reg;
reg [31:0] main_for_cond84_preheader_5;
reg [31:0] main_for_cond84_preheader_5_reg;
reg [31:0] main_for_body86_6;
reg [31:0] main_for_body86_6_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body86_arrayidx88;
reg [31:0] main_for_body86_7;
reg  main_for_body86_cmp89;
reg [31:0] main_for_inc93_8;
reg  main_for_inc93_exitcond67;
reg [6:0] main_for_inc96_9;
reg  main_for_inc96_exitcond69;
reg [5:0] main_for_body101_i_0338;
reg [5:0] main_for_body101_i_0338_reg;
reg [29:0] main_for_body101_bit_select15;
reg [26:0] main_for_body101_bit_select13;
reg [31:0] main_for_body101_bit_concat16;
reg [31:0] main_for_body101_bit_concat14;
reg [31:0] main_for_body101_sr_add;
reg [31:0] main_for_body101_sr_add_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body101_arrayidx102;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body101_arrayidx103;
reg [31:0] main_for_body106_j_0337;
reg [31:0] main_for_body106_j_0337_reg;
reg [31:0] main_for_body106_10;
reg [31:0] main_for_body106_10_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body106_scevgep43;
reg [31:0] main_for_body106_11;
reg [31:0] main_for_body106_11_reg;
reg  main_for_body106_exitcond61;
reg  main_for_body106_exitcond61_reg;
reg [6:0] main_for_inc112_12;
reg  main_for_inc112_exitcond63;
reg [2:0] main_for_cond118_preheader_13;
reg [2:0] main_for_cond118_preheader_13_reg;
reg [26:0] main_for_cond118_preheader_bit_select9;
reg [25:0] main_for_cond118_preheader_bit_select7;
reg [24:0] main_for_cond118_preheader_bit_select5;
reg [3:0] main_for_cond118_preheader_sr_negate;
reg [30:0] main_for_cond118_preheader_bit_select11;
reg [31:0] main_for_cond118_preheader_bit_concat12;
reg [31:0] main_for_cond118_preheader_bit_concat10;
reg [31:0] main_for_cond118_preheader_bit_concat8;
reg [31:0] main_for_cond118_preheader_bit_concat6;
reg [31:0] main_for_cond118_preheader_sr_add82;
reg [31:0] main_for_cond118_preheader_sr_add82_reg;
reg [31:0] main_for_cond118_preheader_sr_add83;
reg [31:0] main_for_cond118_preheader_sr_add83_reg;
reg [31:0] main_for_cond118_preheader_sr_add84;
reg [31:0] main_for_cond118_preheader_sr_add84_reg;
reg [30:0] main_for_cond118_preheader_bit_select3;
reg [31:0] main_for_cond118_preheader_14;
reg [31:0] main_for_cond118_preheader_14_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep41;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep41_reg;
reg [31:0] main_for_cond118_preheader_15;
reg [31:0] main_for_cond118_preheader_15_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep39;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep39_reg;
reg [31:0] main_for_cond118_preheader_16;
reg [31:0] main_for_cond118_preheader_16_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep37;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep37_reg;
reg [31:0] main_for_cond118_preheader_17;
reg [31:0] main_for_cond118_preheader_17_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep36;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep36_reg;
reg [31:0] main_for_cond118_preheader_18;
reg [31:0] main_for_cond118_preheader_18_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep35;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep35_reg;
reg [31:0] main_for_cond118_preheader_19;
reg [31:0] main_for_cond118_preheader_19_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep34;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep34_reg;
reg [31:0] main_for_cond118_preheader_20;
reg [31:0] main_for_cond118_preheader_20_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep33;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep33_reg;
reg [31:0] main_for_cond118_preheader_21;
reg [31:0] main_for_cond118_preheader_21_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep32;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep32_reg;
reg [31:0] main_for_cond118_preheader_22;
reg [31:0] main_for_cond118_preheader_22_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep31;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep31_reg;
reg [31:0] main_for_cond118_preheader_bit_concat4;
reg [31:0] main_for_cond118_preheader_bit_concat4_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond118_preheader_scevgep40;
reg  main_for_cond118_preheader_cmp121;
reg  main_for_cond118_preheader_cmp121_reg;
reg [3:0] main_for_inc192_23;
reg  main_for_inc192_exitcond15;
reg [5:0] main_for_body198_i_2333;
reg [5:0] main_for_body198_i_2333_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body198_arrayidx199;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body198_arrayidx200;
reg [6:0] main_for_body198_inc239;
reg [6:0] main_for_body198_inc239_reg;
reg [31:0] main_for_body198_24;
reg [31:0] main_for_body198_24_reg;
reg [31:0] main_for_body198_25;
reg [31:0] main_for_body198_25_reg;
reg [31:0] main_for_body_i_i_057_i;
reg [31:0] main_for_body_i_i_057_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx1_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_arrayidx2_i;
reg [31:0] main_for_body_i_26;
reg [31:0] main_for_body_i_26_reg;
reg  main_for_body_i_exitcond2;
reg  main_for_body_i_exitcond2_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_end_i_arrayidx_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_end_i_arrayidx3_i;
reg [31:0] main_for_body6_i_count_056_i;
reg [31:0] main_for_body6_i_count_056_i_reg;
reg [31:0] main_for_body_i_i_27;
reg [31:0] main_for_body_i_i_27_reg;
reg [31:0] main_for_body_i_i_min_index_012_i_i;
reg [31:0] main_for_body_i_i_min_index_012_i_i_reg;
reg [31:0] main_for_body_i_i_min_011_i_i;
reg [31:0] main_for_body_i_i_min_011_i_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_i_arrayidx_i_i;
reg [31:0] main_for_body_i_i_28;
reg  main_for_body_i_i_cmp1_i_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_land_lhs_true_i_i_arrayidx2_i_i;
reg [31:0] main_land_lhs_true_i_i_29;
reg  main_land_lhs_true_i_i_cmp3_i_i;
reg [31:0] main_land_lhs_true_i_i_min_0_i_i;
reg [31:0] main_land_lhs_true_i_i_min_index_0_v_0_i_i;
reg [31:0] main_for_inc_i_i_min_1_i_i;
reg [31:0] main_for_inc_i_i_min_1_i_i_reg;
reg [31:0] main_for_inc_i_i_min_index_1_i_i;
reg [31:0] main_for_inc_i_i_min_index_1_i_i_reg;
reg [29:0] main_for_inc_i_i_bit_select1;
reg [29:0] main_for_inc_i_i_bit_select1_reg;
reg [26:0] main_for_inc_i_i_bit_select;
reg [26:0] main_for_inc_i_i_bit_select_reg;
reg [31:0] main_for_inc_i_i_30;
reg  main_for_inc_i_i_exitcond5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_minDistance_exit_i_arrayidx8_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_minDistance_exit_i_arrayidx17_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_minDistance_exit_i_arrayidx17_i_reg;
reg [31:0] main_minDistance_exit_i_bit_concat2;
reg [31:0] main_minDistance_exit_i_bit_concat;
reg [31:0] main_minDistance_exit_i_sr_add87;
reg [31:0] main_minDistance_exit_i_sr_add87_reg;
reg [31:0] main_for_body11_i_v_055_i;
reg [31:0] main_for_body11_i_v_055_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx12_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx20_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx20_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx22_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx22_i_reg;
reg [31:0] main_for_body11_i_31;
reg  main_for_body11_i_tobool_i;
reg [31:0] main_land_lhs_true_i_32;
reg [31:0] main_land_lhs_true_i_32_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_land_lhs_true_i_scevgep;
reg [31:0] main_land_lhs_true_i_33;
reg [31:0] main_land_lhs_true_i_33_reg;
reg  main_land_lhs_true_i_tobool15_i;
reg [31:0] main_land_lhs_true16_i_34;
reg [31:0] main_land_lhs_true16_i_add_i;
reg [31:0] main_land_lhs_true16_i_add_i_reg;
reg [31:0] main_land_lhs_true16_i_35;
reg  main_land_lhs_true16_i_cmp21_i;
reg [31:0] main_for_inc28_i_36;
reg  main_for_inc28_i_exitcond8;
reg [31:0] main_for_inc31_i_37;
reg  main_for_inc31_i_exitcond;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_dijkstra_exit_arrayidx207329;
reg [31:0] main_dijkstra_exit_38;
reg [31:0] main_dijkstra_exit_38_reg;
reg  main_dijkstra_exit_cmp208330;
reg [31:0] main_if_end211_39;
reg [31:0] main_if_end211_39_reg;
reg [31:0] main_if_end211_origem_1332;
reg [31:0] main_if_end211_origem_1332_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end211_arrayidx212;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end211_arrayidx212_reg;
reg [31:0] main_if_end211_40;
reg [31:0] main_if_end211_40_reg;
reg  main_if_end211_cmp213;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end211_arrayidx215;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end211_arrayidx215_reg;
reg [31:0] main_if_end211_41;
reg [31:0] main_if_end211_41_reg;
reg  main_if_end211_cmp216;
reg  main_if_end211_and218323;
reg [31:0] main_if_then220_add228;
reg [31:0] main_if_then220_add230;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then220_arrayidx207;
reg [31:0] main_if_then220_42;
reg  main_if_then220_cmp208;
reg  main_for_inc238_cmp196;
reg [31:0] main_for_inc189_us_5_43;
reg [31:0] main_for_inc189_us_5_43_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep38;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep38_reg;
reg [31:0] main_for_inc189_us_5_44;
reg [31:0] main_for_inc189_us_5_44_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep30;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep30_reg;
reg [31:0] main_for_inc189_us_5_45;
reg [31:0] main_for_inc189_us_5_45_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep29;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep29_reg;
reg [31:0] main_for_inc189_us_5_46;
reg [31:0] main_for_inc189_us_5_46_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep28;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep28_reg;
reg [31:0] main_for_inc189_us_5_47;
reg [31:0] main_for_inc189_us_5_47_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep27;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep27_reg;
reg [31:0] main_for_inc189_us_5_48;
reg [31:0] main_for_inc189_us_5_48_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep26;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep26_reg;
reg [31:0] main_for_inc189_us_5_49;
reg [31:0] main_for_inc189_us_5_49_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep25;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep25_reg;
reg [31:0] main_for_inc189_us_5_50;
reg [31:0] main_for_inc189_us_5_50_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep24;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep24_reg;
reg [31:0] main_for_inc189_us_5_51;
reg [31:0] main_for_inc189_us_5_51_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep23;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep23_reg;
reg [31:0] main_for_inc189_us_5_52;
reg [31:0] main_for_inc189_us_5_52_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep22;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep22_reg;
reg [31:0] main_for_inc189_us_5_53;
reg [31:0] main_for_inc189_us_5_53_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep21;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep21_reg;
reg [31:0] main_for_inc189_us_5_54;
reg [31:0] main_for_inc189_us_5_54_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep20;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc189_us_5_scevgep20_reg;
reg [5:0] main_grid_address_a;
wire [31:0] main_grid_out_a;
wire [5:0] main_grid_address_b;
wire [31:0] main_grid_out_b;
reg [5:0] main_entry_dist_i_address_a;
reg  main_entry_dist_i_write_enable_a;
reg [31:0] main_entry_dist_i_in_a;
wire [31:0] main_entry_dist_i_out_a;
reg [5:0] main_entry_dist_i_address_b;
reg  main_entry_dist_i_write_enable_b;
reg [31:0] main_entry_dist_i_in_b;
wire [31:0] main_entry_dist_i_out_b;
reg [5:0] main_entry_sptSet_i_address_a;
reg  main_entry_sptSet_i_write_enable_a;
reg [31:0] main_entry_sptSet_i_in_a;
wire [31:0] main_entry_sptSet_i_out_a;
reg [5:0] main_entry_parent_address_a;
reg  main_entry_parent_write_enable_a;
reg [31:0] main_entry_parent_in_a;
wire [31:0] main_entry_parent_out_a;
reg [10:0] main_entry_m1_address_a;
reg  main_entry_m1_write_enable_a;
reg [31:0] main_entry_m1_in_a;
wire [31:0] main_entry_m1_out_a;
reg [10:0] main_entry_m1_address_b;
reg  main_entry_m1_write_enable_b;
reg [31:0] main_entry_m1_in_b;
wire [31:0] main_entry_m1_out_b;
reg [5:0] main_entry_indice_e_address_a;
reg  main_entry_indice_e_write_enable_a;
reg [31:0] main_entry_indice_e_in_a;
wire [31:0] main_entry_indice_e_out_a;
reg [5:0] main_entry_indice_s_address_a;
reg  main_entry_indice_s_write_enable_a;
reg [31:0] main_entry_indice_s_in_a;
wire [31:0] main_entry_indice_s_out_a;
reg [4:0] main_entry_vla319_address_a;
reg  main_entry_vla319_write_enable_a;
reg [31:0] main_entry_vla319_in_a;
wire [31:0] main_entry_vla319_out_a;
reg [4:0] main_entry_vla319_address_b;
reg  main_entry_vla319_write_enable_b;
reg [31:0] main_entry_vla319_in_b;
wire [31:0] main_entry_vla319_out_b;
reg [4:0] main_entry_vla1320_address_a;
reg  main_entry_vla1320_write_enable_a;
reg [31:0] main_entry_vla1320_in_a;
wire [31:0] main_entry_vla1320_out_a;
reg [4:0] main_entry_vla1320_address_b;
reg  main_entry_vla1320_write_enable_b;
reg [31:0] main_entry_vla1320_in_b;
wire [31:0] main_entry_vla1320_out_b;
reg [4:0] main_entry_vla65321_address_a;
reg  main_entry_vla65321_write_enable_a;
reg [31:0] main_entry_vla65321_in_a;
wire [31:0] main_entry_vla65321_out_a;
reg [4:0] main_entry_vla66322_address_a;
reg  main_entry_vla66322_write_enable_a;
reg [31:0] main_entry_vla66322_in_a;
wire [31:0] main_entry_vla66322_out_a;
reg [29:0] main_for_body101_i_0338_reg_width_extended;
wire [1:0] main_for_body101_bit_concat16_bit_select_operand_2;
wire [4:0] main_for_body101_bit_concat14_bit_select_operand_2;
reg [26:0] main_for_cond118_preheader_13_reg_width_extended;
reg [30:0] main_for_cond118_preheader_sr_negate_width_extended;
wire  main_for_cond118_preheader_bit_concat12_bit_select_operand_2;
wire [4:0] main_for_cond118_preheader_bit_concat10_bit_select_operand_2;
wire [5:0] main_for_cond118_preheader_bit_concat8_bit_select_operand_2;
wire [6:0] main_for_cond118_preheader_bit_concat6_bit_select_operand_2;
reg [3:0] main_for_cond118_preheader_cmp121_op0_temp;
wire [4:0] main_for_cond118_preheader_cmp121_op1_temp;
wire  main_for_cond118_preheader_bit_concat4_bit_select_operand_2;
wire [1:0] main_minDistance_exit_i_bit_concat2_bit_select_operand_2;
wire [4:0] main_minDistance_exit_i_bit_concat_bit_select_operand_2;
wire [4:0] main_if_end211_cmp213_op1_temp;
wire [4:0] main_if_end211_cmp216_op1_temp;
reg [7:0] main_for_inc238_cmp196_op0_temp;
wire [7:0] main_for_inc238_cmp196_op1_temp;



// @main.grid = private unnamed_addr constant [36 x i32] [i32 21, i32 23, i32 7, i32 20, i32 15, i32 13, i32 26, i32 25, i32 24, i32 18, i32 9, i32 5, i32 16, i32 17, i32 2, i32 11, i32 1, i32 3, i32 255...
rom_dual_port main_grid (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_grid_address_a ),
	.q_a( main_grid_out_a ),
	.address_b( main_grid_address_b ),
	.q_b( main_grid_out_b )
);
defparam main_grid.width_a = 32;
defparam main_grid.widthad_a = 6;
defparam main_grid.numwords_a = 36;
defparam main_grid.width_b = 32;
defparam main_grid.widthad_b = 6;
defparam main_grid.numwords_b = 36;
defparam main_grid.latency = 1;
defparam main_grid.init_file = {`MEM_INIT_DIR, "main_grid.mif"};


//   %dist.i = alloca [36 x i32], align 4, !dbg !83, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_dist_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_dist_i_address_a ),
	.wren_a( main_entry_dist_i_write_enable_a ),
	.data_a( main_entry_dist_i_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_dist_i_out_a ),
	.address_b( main_entry_dist_i_address_b ),
	.wren_b( main_entry_dist_i_write_enable_b ),
	.data_b( main_entry_dist_i_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_dist_i_out_b )
);
defparam main_entry_dist_i.width_a = 32;
defparam main_entry_dist_i.widthad_a = 6;
defparam main_entry_dist_i.width_be_a = 4;
defparam main_entry_dist_i.numwords_a = 36;
defparam main_entry_dist_i.width_b = 32;
defparam main_entry_dist_i.widthad_b = 6;
defparam main_entry_dist_i.width_be_b = 4;
defparam main_entry_dist_i.numwords_b = 36;
defparam main_entry_dist_i.latency = 1;


//   %sptSet.i = alloca [36 x i32], align 4, !dbg !83, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_sptSet_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_sptSet_i_address_a ),
	.wren_a( main_entry_sptSet_i_write_enable_a ),
	.data_a( main_entry_sptSet_i_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_sptSet_i_out_a )
);
defparam main_entry_sptSet_i.width_a = 32;
defparam main_entry_sptSet_i.widthad_a = 6;
defparam main_entry_sptSet_i.width_be_a = 4;
defparam main_entry_sptSet_i.numwords_a = 36;
defparam main_entry_sptSet_i.latency = 1;


//   %parent = alloca [36 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_parent (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_parent_address_a ),
	.wren_a( main_entry_parent_write_enable_a ),
	.data_a( main_entry_parent_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_parent_out_a )
);
defparam main_entry_parent.width_a = 32;
defparam main_entry_parent.widthad_a = 6;
defparam main_entry_parent.width_be_a = 4;
defparam main_entry_parent.numwords_a = 36;
defparam main_entry_parent.latency = 1;


//   %m1 = alloca [1296 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_m1 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_m1_address_a ),
	.wren_a( main_entry_m1_write_enable_a ),
	.data_a( main_entry_m1_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_m1_out_a ),
	.address_b( main_entry_m1_address_b ),
	.wren_b( main_entry_m1_write_enable_b ),
	.data_b( main_entry_m1_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_m1_out_b )
);
defparam main_entry_m1.width_a = 32;
defparam main_entry_m1.widthad_a = 11;
defparam main_entry_m1.width_be_a = 4;
defparam main_entry_m1.numwords_a = 1296;
defparam main_entry_m1.width_b = 32;
defparam main_entry_m1.widthad_b = 11;
defparam main_entry_m1.width_be_b = 4;
defparam main_entry_m1.numwords_b = 1296;
defparam main_entry_m1.latency = 1;


//   %indice_e = alloca [36 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_indice_e (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_indice_e_address_a ),
	.wren_a( main_entry_indice_e_write_enable_a ),
	.data_a( main_entry_indice_e_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_indice_e_out_a )
);
defparam main_entry_indice_e.width_a = 32;
defparam main_entry_indice_e.widthad_a = 6;
defparam main_entry_indice_e.width_be_a = 4;
defparam main_entry_indice_e.numwords_a = 36;
defparam main_entry_indice_e.latency = 1;


//   %indice_s = alloca [36 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_indice_s (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_indice_s_address_a ),
	.wren_a( main_entry_indice_s_write_enable_a ),
	.data_a( main_entry_indice_s_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_indice_s_out_a )
);
defparam main_entry_indice_s.width_a = 32;
defparam main_entry_indice_s.widthad_a = 6;
defparam main_entry_indice_s.width_be_a = 4;
defparam main_entry_indice_s.numwords_a = 36;
defparam main_entry_indice_s.latency = 1;


//   %vla319 = alloca [32 x i32], align 4, !dbg !88, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_vla319 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla319_address_a ),
	.wren_a( main_entry_vla319_write_enable_a ),
	.data_a( main_entry_vla319_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla319_out_a ),
	.address_b( main_entry_vla319_address_b ),
	.wren_b( main_entry_vla319_write_enable_b ),
	.data_b( main_entry_vla319_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_vla319_out_b )
);
defparam main_entry_vla319.width_a = 32;
defparam main_entry_vla319.widthad_a = 5;
defparam main_entry_vla319.width_be_a = 4;
defparam main_entry_vla319.numwords_a = 32;
defparam main_entry_vla319.width_b = 32;
defparam main_entry_vla319.widthad_b = 5;
defparam main_entry_vla319.width_be_b = 4;
defparam main_entry_vla319.numwords_b = 32;
defparam main_entry_vla319.latency = 1;


//   %vla1320 = alloca [32 x i32], align 4, !dbg !89, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_vla1320 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla1320_address_a ),
	.wren_a( main_entry_vla1320_write_enable_a ),
	.data_a( main_entry_vla1320_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla1320_out_a ),
	.address_b( main_entry_vla1320_address_b ),
	.wren_b( main_entry_vla1320_write_enable_b ),
	.data_b( main_entry_vla1320_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_vla1320_out_b )
);
defparam main_entry_vla1320.width_a = 32;
defparam main_entry_vla1320.widthad_a = 5;
defparam main_entry_vla1320.width_be_a = 4;
defparam main_entry_vla1320.numwords_a = 32;
defparam main_entry_vla1320.width_b = 32;
defparam main_entry_vla1320.widthad_b = 5;
defparam main_entry_vla1320.width_be_b = 4;
defparam main_entry_vla1320.numwords_b = 32;
defparam main_entry_vla1320.latency = 1;


//   %vla65321 = alloca [32 x i32], align 4, !dbg !158, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_vla65321 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla65321_address_a ),
	.wren_a( main_entry_vla65321_write_enable_a ),
	.data_a( main_entry_vla65321_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla65321_out_a )
);
defparam main_entry_vla65321.width_a = 32;
defparam main_entry_vla65321.widthad_a = 5;
defparam main_entry_vla65321.width_be_a = 4;
defparam main_entry_vla65321.numwords_a = 32;
defparam main_entry_vla65321.latency = 1;


//   %vla66322 = alloca [32 x i32], align 4, !dbg !158, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_vla66322 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla66322_address_a ),
	.wren_a( main_entry_vla66322_write_enable_a ),
	.data_a( main_entry_vla66322_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla66322_out_a )
);
defparam main_entry_vla66322.width_a = 32;
defparam main_entry_vla66322.widthad_a = 5;
defparam main_entry_vla66322.width_be_a = 4;
defparam main_entry_vla66322.numwords_a = 32;
defparam main_entry_vla66322.latency = 1;

always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_entry_1;
LEGUP_F_main_BB_dijkstra_exit_75:
		next_state = LEGUP_F_main_BB_dijkstra_exit_76;
LEGUP_F_main_BB_dijkstra_exit_76:
	if ((fsm_stall == 1'd0) && (main_dijkstra_exit_cmp208330 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc238_83;
	else if ((fsm_stall == 1'd0) && (main_dijkstra_exit_cmp208330 == 1'd0))
		next_state = LEGUP_F_main_BB_if_end211_preheader_77;
LEGUP_F_main_BB_entry_1:
		next_state = LEGUP_F_main_BB_entry_2;
LEGUP_F_main_BB_entry_10:
		next_state = LEGUP_F_main_BB_entry_11;
LEGUP_F_main_BB_entry_11:
		next_state = LEGUP_F_main_BB_entry_12;
LEGUP_F_main_BB_entry_12:
		next_state = LEGUP_F_main_BB_entry_13;
LEGUP_F_main_BB_entry_13:
		next_state = LEGUP_F_main_BB_entry_14;
LEGUP_F_main_BB_entry_14:
		next_state = LEGUP_F_main_BB_entry_15;
LEGUP_F_main_BB_entry_15:
		next_state = LEGUP_F_main_BB_entry_16;
LEGUP_F_main_BB_entry_16:
		next_state = LEGUP_F_main_BB_entry_17;
LEGUP_F_main_BB_entry_17:
		next_state = LEGUP_F_main_BB_for_cond69_preheader_18;
LEGUP_F_main_BB_entry_2:
		next_state = LEGUP_F_main_BB_entry_3;
LEGUP_F_main_BB_entry_3:
		next_state = LEGUP_F_main_BB_entry_4;
LEGUP_F_main_BB_entry_4:
		next_state = LEGUP_F_main_BB_entry_5;
LEGUP_F_main_BB_entry_5:
		next_state = LEGUP_F_main_BB_entry_6;
LEGUP_F_main_BB_entry_6:
		next_state = LEGUP_F_main_BB_entry_7;
LEGUP_F_main_BB_entry_7:
		next_state = LEGUP_F_main_BB_entry_8;
LEGUP_F_main_BB_entry_8:
		next_state = LEGUP_F_main_BB_entry_9;
LEGUP_F_main_BB_entry_9:
		next_state = LEGUP_F_main_BB_entry_10;
LEGUP_F_main_BB_for_body101_36:
		next_state = LEGUP_F_main_BB_for_body101_37;
LEGUP_F_main_BB_for_body101_37:
		next_state = LEGUP_F_main_BB_for_body106_38;
LEGUP_F_main_BB_for_body101_preheader_35:
		next_state = LEGUP_F_main_BB_for_body101_36;
LEGUP_F_main_BB_for_body106_38:
		next_state = LEGUP_F_main_BB_for_body106_39;
LEGUP_F_main_BB_for_body106_39:
		next_state = LEGUP_F_main_BB_for_body106_40;
LEGUP_F_main_BB_for_body106_40:
	if ((fsm_stall == 1'd0) && (main_for_body106_exitcond61_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc112_41;
	else if ((fsm_stall == 1'd0) && (main_for_body106_exitcond61_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body106_38;
LEGUP_F_main_BB_for_body11_i_64:
		next_state = LEGUP_F_main_BB_for_body11_i_65;
LEGUP_F_main_BB_for_body11_i_65:
	if ((fsm_stall == 1'd0) && (main_for_body11_i_tobool_i == 1'd1))
		next_state = LEGUP_F_main_BB_land_lhs_true_i_66;
	else if ((fsm_stall == 1'd0) && (main_for_body11_i_tobool_i == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc28_i_73;
LEGUP_F_main_BB_for_body198_50:
		next_state = LEGUP_F_main_BB_for_body198_51;
LEGUP_F_main_BB_for_body198_51:
		next_state = LEGUP_F_main_BB_for_body_i_52;
LEGUP_F_main_BB_for_body198_preheader_49:
		next_state = LEGUP_F_main_BB_for_body198_50;
LEGUP_F_main_BB_for_body6_i_56:
		next_state = LEGUP_F_main_BB_for_body_i_i_57;
LEGUP_F_main_BB_for_body71_20:
		next_state = LEGUP_F_main_BB_for_body71_21;
LEGUP_F_main_BB_for_body71_21:
	if ((fsm_stall == 1'd0) && (main_for_body71_cmp74 == 1'd1))
		next_state = LEGUP_F_main_BB_if_then_22;
	else if ((fsm_stall == 1'd0) && (main_for_body71_cmp74 == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc_24;
LEGUP_F_main_BB_for_body86_29:
		next_state = LEGUP_F_main_BB_for_body86_30;
LEGUP_F_main_BB_for_body86_30:
	if ((fsm_stall == 1'd0) && (main_for_body86_cmp89 == 1'd1))
		next_state = LEGUP_F_main_BB_if_then90_31;
	else if ((fsm_stall == 1'd0) && (main_for_body86_cmp89 == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc93_33;
LEGUP_F_main_BB_for_body_i_52:
		next_state = LEGUP_F_main_BB_for_body_i_53;
LEGUP_F_main_BB_for_body_i_53:
	if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond2_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_end_i_54;
	else if ((fsm_stall == 1'd0) && (main_for_body_i_exitcond2_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_i_52;
LEGUP_F_main_BB_for_body_i_i_57:
		next_state = LEGUP_F_main_BB_for_body_i_i_58;
LEGUP_F_main_BB_for_body_i_i_58:
	if ((fsm_stall == 1'd0) && (main_for_body_i_i_cmp1_i_i == 1'd1))
		next_state = LEGUP_F_main_BB_land_lhs_true_i_i_59;
	else if ((fsm_stall == 1'd0) && (main_for_body_i_i_cmp1_i_i == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc_i_i_61;
LEGUP_F_main_BB_for_cond118_preheader_43:
		next_state = LEGUP_F_main_BB_for_cond118_preheader_44;
LEGUP_F_main_BB_for_cond118_preheader_44:
		next_state = LEGUP_F_main_BB_for_cond118_preheader_45;
LEGUP_F_main_BB_for_cond118_preheader_45:
		next_state = LEGUP_F_main_BB_for_cond118_preheader_46;
LEGUP_F_main_BB_for_cond118_preheader_46:
		next_state = LEGUP_F_main_BB_for_cond118_preheader_47;
LEGUP_F_main_BB_for_cond118_preheader_47:
	if ((fsm_stall == 1'd0) && (main_for_cond118_preheader_cmp121_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc189_us_5_92;
	else if ((fsm_stall == 1'd0) && (main_for_cond118_preheader_cmp121_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc189_5_87;
LEGUP_F_main_BB_for_cond118_preheader_preheader_42:
		next_state = LEGUP_F_main_BB_for_cond118_preheader_43;
LEGUP_F_main_BB_for_cond69_preheader_18:
		next_state = LEGUP_F_main_BB_for_cond69_preheader_19;
LEGUP_F_main_BB_for_cond69_preheader_19:
		next_state = LEGUP_F_main_BB_for_body71_20;
LEGUP_F_main_BB_for_cond84_preheader_27:
		next_state = LEGUP_F_main_BB_for_cond84_preheader_28;
LEGUP_F_main_BB_for_cond84_preheader_28:
		next_state = LEGUP_F_main_BB_for_body86_29;
LEGUP_F_main_BB_for_cond84_preheader_preheader_26:
		next_state = LEGUP_F_main_BB_for_cond84_preheader_27;
LEGUP_F_main_BB_for_end240_86:
		next_state = LEGUP_0;
LEGUP_F_main_BB_for_end240_loopexit1_85:
		next_state = LEGUP_F_main_BB_for_end240_86;
LEGUP_F_main_BB_for_end240_loopexit_84:
		next_state = LEGUP_F_main_BB_for_end240_86;
LEGUP_F_main_BB_for_end_i_54:
		next_state = LEGUP_F_main_BB_for_end_i_55;
LEGUP_F_main_BB_for_end_i_55:
		next_state = LEGUP_F_main_BB_for_body6_i_56;
LEGUP_F_main_BB_for_inc112_41:
	if ((fsm_stall == 1'd0) && (main_for_inc112_exitcond63 == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond118_preheader_preheader_42;
	else if ((fsm_stall == 1'd0) && (main_for_inc112_exitcond63 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body101_36;
LEGUP_F_main_BB_for_inc189_5_87:
		next_state = LEGUP_F_main_BB_for_inc189_5_88;
LEGUP_F_main_BB_for_inc189_5_88:
		next_state = LEGUP_F_main_BB_for_inc189_5_89;
LEGUP_F_main_BB_for_inc189_5_89:
		next_state = LEGUP_F_main_BB_for_inc189_5_90;
LEGUP_F_main_BB_for_inc189_5_90:
		next_state = LEGUP_F_main_BB_for_inc189_5_91;
LEGUP_F_main_BB_for_inc189_5_91:
		next_state = LEGUP_F_main_BB_for_inc192_48;
LEGUP_F_main_BB_for_inc189_us_5_100:
		next_state = LEGUP_F_main_BB_for_inc189_us_5_101;
LEGUP_F_main_BB_for_inc189_us_5_101:
		next_state = LEGUP_F_main_BB_for_inc189_us_5_102;
LEGUP_F_main_BB_for_inc189_us_5_102:
		next_state = LEGUP_F_main_BB_for_inc192_48;
LEGUP_F_main_BB_for_inc189_us_5_92:
		next_state = LEGUP_F_main_BB_for_inc189_us_5_93;
LEGUP_F_main_BB_for_inc189_us_5_93:
		next_state = LEGUP_F_main_BB_for_inc189_us_5_94;
LEGUP_F_main_BB_for_inc189_us_5_94:
		next_state = LEGUP_F_main_BB_for_inc189_us_5_95;
LEGUP_F_main_BB_for_inc189_us_5_95:
		next_state = LEGUP_F_main_BB_for_inc189_us_5_96;
LEGUP_F_main_BB_for_inc189_us_5_96:
		next_state = LEGUP_F_main_BB_for_inc189_us_5_97;
LEGUP_F_main_BB_for_inc189_us_5_97:
		next_state = LEGUP_F_main_BB_for_inc189_us_5_98;
LEGUP_F_main_BB_for_inc189_us_5_98:
		next_state = LEGUP_F_main_BB_for_inc189_us_5_99;
LEGUP_F_main_BB_for_inc189_us_5_99:
		next_state = LEGUP_F_main_BB_for_inc189_us_5_100;
LEGUP_F_main_BB_for_inc192_48:
	if ((fsm_stall == 1'd0) && (main_for_inc192_exitcond15 == 1'd1))
		next_state = LEGUP_F_main_BB_for_body198_preheader_49;
	else if ((fsm_stall == 1'd0) && (main_for_inc192_exitcond15 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond118_preheader_43;
LEGUP_F_main_BB_for_inc238_83:
	if ((fsm_stall == 1'd0) && (main_for_inc238_cmp196 == 1'd1))
		next_state = LEGUP_F_main_BB_for_body198_50;
	else if ((fsm_stall == 1'd0) && (main_for_inc238_cmp196 == 1'd0))
		next_state = LEGUP_F_main_BB_for_end240_loopexit1_85;
LEGUP_F_main_BB_for_inc238_loopexit_82:
		next_state = LEGUP_F_main_BB_for_inc238_83;
LEGUP_F_main_BB_for_inc28_i_73:
	if ((fsm_stall == 1'd0) && (main_for_inc28_i_exitcond8 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc31_i_74;
	else if ((fsm_stall == 1'd0) && (main_for_inc28_i_exitcond8 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body11_i_64;
LEGUP_F_main_BB_for_inc31_i_74:
	if ((fsm_stall == 1'd0) && (main_for_inc31_i_exitcond == 1'd1))
		next_state = LEGUP_F_main_BB_dijkstra_exit_75;
	else if ((fsm_stall == 1'd0) && (main_for_inc31_i_exitcond == 1'd0))
		next_state = LEGUP_F_main_BB_for_body6_i_56;
LEGUP_F_main_BB_for_inc76_25:
	if ((fsm_stall == 1'd0) && (main_for_inc76_exitcond74 == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond84_preheader_preheader_26;
	else if ((fsm_stall == 1'd0) && (main_for_inc76_exitcond74 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond69_preheader_18;
LEGUP_F_main_BB_for_inc93_33:
	if ((fsm_stall == 1'd0) && (main_for_inc93_exitcond67 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc96_34;
	else if ((fsm_stall == 1'd0) && (main_for_inc93_exitcond67 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body86_29;
LEGUP_F_main_BB_for_inc96_34:
	if ((fsm_stall == 1'd0) && (main_for_inc96_exitcond69 == 1'd1))
		next_state = LEGUP_F_main_BB_for_body101_preheader_35;
	else if ((fsm_stall == 1'd0) && (main_for_inc96_exitcond69 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond84_preheader_27;
LEGUP_F_main_BB_for_inc_24:
	if ((fsm_stall == 1'd0) && (main_for_inc_exitcond72 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc76_25;
	else if ((fsm_stall == 1'd0) && (main_for_inc_exitcond72 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body71_20;
LEGUP_F_main_BB_for_inc_i_i_61:
	if ((fsm_stall == 1'd0) && (main_for_inc_i_i_exitcond5 == 1'd1))
		next_state = LEGUP_F_main_BB_minDistance_exit_i_62;
	else if ((fsm_stall == 1'd0) && (main_for_inc_i_i_exitcond5 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_i_i_57;
LEGUP_F_main_BB_if_end211_78:
		next_state = LEGUP_F_main_BB_if_end211_79;
LEGUP_F_main_BB_if_end211_79:
	if ((fsm_stall == 1'd0) && (main_if_end211_and218323 == 1'd1))
		next_state = LEGUP_F_main_BB_if_then220_80;
	else if ((fsm_stall == 1'd0) && (main_if_end211_and218323 == 1'd0))
		next_state = LEGUP_F_main_BB_for_end240_loopexit_84;
LEGUP_F_main_BB_if_end211_preheader_77:
		next_state = LEGUP_F_main_BB_if_end211_78;
LEGUP_F_main_BB_if_then220_80:
		next_state = LEGUP_F_main_BB_if_then220_81;
LEGUP_F_main_BB_if_then220_81:
	if ((fsm_stall == 1'd0) && (main_if_then220_cmp208 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc238_loopexit_82;
	else if ((fsm_stall == 1'd0) && (main_if_then220_cmp208 == 1'd0))
		next_state = LEGUP_F_main_BB_if_end211_78;
LEGUP_F_main_BB_if_then90_31:
		next_state = LEGUP_F_main_BB_if_then90_32;
LEGUP_F_main_BB_if_then90_32:
		next_state = LEGUP_F_main_BB_for_inc93_33;
LEGUP_F_main_BB_if_then_22:
		next_state = LEGUP_F_main_BB_if_then_23;
LEGUP_F_main_BB_if_then_23:
		next_state = LEGUP_F_main_BB_for_inc_24;
LEGUP_F_main_BB_if_then_i_71:
		next_state = LEGUP_F_main_BB_if_then_i_72;
LEGUP_F_main_BB_if_then_i_72:
		next_state = LEGUP_F_main_BB_for_inc28_i_73;
LEGUP_F_main_BB_land_lhs_true16_i_69:
		next_state = LEGUP_F_main_BB_land_lhs_true16_i_70;
LEGUP_F_main_BB_land_lhs_true16_i_70:
	if ((fsm_stall == 1'd0) && (main_land_lhs_true16_i_cmp21_i == 1'd1))
		next_state = LEGUP_F_main_BB_if_then_i_71;
	else if ((fsm_stall == 1'd0) && (main_land_lhs_true16_i_cmp21_i == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc28_i_73;
LEGUP_F_main_BB_land_lhs_true_i_66:
		next_state = LEGUP_F_main_BB_land_lhs_true_i_67;
LEGUP_F_main_BB_land_lhs_true_i_67:
		next_state = LEGUP_F_main_BB_land_lhs_true_i_68;
LEGUP_F_main_BB_land_lhs_true_i_68:
	if ((fsm_stall == 1'd0) && (main_land_lhs_true_i_tobool15_i == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc28_i_73;
	else if ((fsm_stall == 1'd0) && (main_land_lhs_true_i_tobool15_i == 1'd0))
		next_state = LEGUP_F_main_BB_land_lhs_true16_i_69;
LEGUP_F_main_BB_land_lhs_true_i_i_59:
		next_state = LEGUP_F_main_BB_land_lhs_true_i_i_60;
LEGUP_F_main_BB_land_lhs_true_i_i_60:
		next_state = LEGUP_F_main_BB_for_inc_i_i_61;
LEGUP_F_main_BB_minDistance_exit_i_62:
		next_state = LEGUP_F_main_BB_minDistance_exit_i_63;
LEGUP_F_main_BB_minDistance_exit_i_63:
		next_state = LEGUP_F_main_BB_for_body11_i_64;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
assign main_entry_vla1320_sub = 1'd0;
assign main_entry_vla319_sub = 1'd0;
assign main_entry_arrayidx3 = (1'd0 + (4 * 32'd1));
assign main_entry_arrayidx4 = (1'd0 + (4 * 32'd1));
assign main_entry_arrayidx5 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx5_reg <= main_entry_arrayidx5;
	end
end
assign main_entry_arrayidx6 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx6_reg <= main_entry_arrayidx6;
	end
end
assign main_entry_arrayidx7 = (1'd0 + (4 * 32'd3));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx7_reg <= main_entry_arrayidx7;
	end
end
assign main_entry_arrayidx8 = (1'd0 + (4 * 32'd3));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx8_reg <= main_entry_arrayidx8;
	end
end
assign main_entry_arrayidx9 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx9_reg <= main_entry_arrayidx9;
	end
end
assign main_entry_arrayidx10 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx10_reg <= main_entry_arrayidx10;
	end
end
assign main_entry_arrayidx11 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx11_reg <= main_entry_arrayidx11;
	end
end
assign main_entry_arrayidx12 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx12_reg <= main_entry_arrayidx12;
	end
end
assign main_entry_arrayidx13 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx13_reg <= main_entry_arrayidx13;
	end
end
assign main_entry_arrayidx14 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx14_reg <= main_entry_arrayidx14;
	end
end
assign main_entry_arrayidx15 = (1'd0 + (4 * 32'd7));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx15_reg <= main_entry_arrayidx15;
	end
end
assign main_entry_arrayidx16 = (1'd0 + (4 * 32'd7));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx16_reg <= main_entry_arrayidx16;
	end
end
assign main_entry_arrayidx17 = (1'd0 + (4 * 32'd8));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx17_reg <= main_entry_arrayidx17;
	end
end
assign main_entry_arrayidx18 = (1'd0 + (4 * 32'd8));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx18_reg <= main_entry_arrayidx18;
	end
end
assign main_entry_arrayidx19 = (1'd0 + (4 * 32'd9));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx19_reg <= main_entry_arrayidx19;
	end
end
assign main_entry_arrayidx20 = (1'd0 + (4 * 32'd9));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx20_reg <= main_entry_arrayidx20;
	end
end
assign main_entry_arrayidx21 = (1'd0 + (4 * 32'd10));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx21_reg <= main_entry_arrayidx21;
	end
end
assign main_entry_arrayidx22 = (1'd0 + (4 * 32'd10));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx22_reg <= main_entry_arrayidx22;
	end
end
assign main_entry_arrayidx23 = (1'd0 + (4 * 32'd11));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx23_reg <= main_entry_arrayidx23;
	end
end
assign main_entry_arrayidx24 = (1'd0 + (4 * 32'd11));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx24_reg <= main_entry_arrayidx24;
	end
end
assign main_entry_arrayidx25 = (1'd0 + (4 * 32'd12));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx25_reg <= main_entry_arrayidx25;
	end
end
assign main_entry_arrayidx26 = (1'd0 + (4 * 32'd12));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx26_reg <= main_entry_arrayidx26;
	end
end
assign main_entry_arrayidx27 = (1'd0 + (4 * 32'd13));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx27_reg <= main_entry_arrayidx27;
	end
end
assign main_entry_arrayidx28 = (1'd0 + (4 * 32'd13));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx28_reg <= main_entry_arrayidx28;
	end
end
assign main_entry_arrayidx29 = (1'd0 + (4 * 32'd14));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx29_reg <= main_entry_arrayidx29;
	end
end
assign main_entry_arrayidx30 = (1'd0 + (4 * 32'd14));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx30_reg <= main_entry_arrayidx30;
	end
end
assign main_entry_arrayidx31 = (1'd0 + (4 * 32'd15));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx31_reg <= main_entry_arrayidx31;
	end
end
assign main_entry_arrayidx32 = (1'd0 + (4 * 32'd15));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx32_reg <= main_entry_arrayidx32;
	end
end
assign main_entry_arrayidx33 = (1'd0 + (4 * 32'd16));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx33_reg <= main_entry_arrayidx33;
	end
end
assign main_entry_arrayidx34 = (1'd0 + (4 * 32'd16));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx34_reg <= main_entry_arrayidx34;
	end
end
assign main_entry_arrayidx35 = (1'd0 + (4 * 32'd17));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx35_reg <= main_entry_arrayidx35;
	end
end
assign main_entry_arrayidx36 = (1'd0 + (4 * 32'd17));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx36_reg <= main_entry_arrayidx36;
	end
end
assign main_entry_arrayidx37 = (1'd0 + (4 * 32'd18));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx37_reg <= main_entry_arrayidx37;
	end
end
assign main_entry_arrayidx38 = (1'd0 + (4 * 32'd18));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx38_reg <= main_entry_arrayidx38;
	end
end
assign main_entry_arrayidx39 = (1'd0 + (4 * 32'd19));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx39_reg <= main_entry_arrayidx39;
	end
end
assign main_entry_arrayidx40 = (1'd0 + (4 * 32'd19));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx40_reg <= main_entry_arrayidx40;
	end
end
assign main_entry_arrayidx41 = (1'd0 + (4 * 32'd20));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx41_reg <= main_entry_arrayidx41;
	end
end
assign main_entry_arrayidx42 = (1'd0 + (4 * 32'd20));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx42_reg <= main_entry_arrayidx42;
	end
end
assign main_entry_arrayidx43 = (1'd0 + (4 * 32'd21));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx43_reg <= main_entry_arrayidx43;
	end
end
assign main_entry_arrayidx44 = (1'd0 + (4 * 32'd21));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx44_reg <= main_entry_arrayidx44;
	end
end
assign main_entry_arrayidx45 = (1'd0 + (4 * 32'd22));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx45_reg <= main_entry_arrayidx45;
	end
end
assign main_entry_arrayidx46 = (1'd0 + (4 * 32'd22));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx46_reg <= main_entry_arrayidx46;
	end
end
assign main_entry_arrayidx47 = (1'd0 + (4 * 32'd23));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx47_reg <= main_entry_arrayidx47;
	end
end
assign main_entry_arrayidx48 = (1'd0 + (4 * 32'd23));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx48_reg <= main_entry_arrayidx48;
	end
end
assign main_entry_arrayidx49 = (1'd0 + (4 * 32'd24));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx49_reg <= main_entry_arrayidx49;
	end
end
assign main_entry_arrayidx50 = (1'd0 + (4 * 32'd24));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx50_reg <= main_entry_arrayidx50;
	end
end
assign main_entry_arrayidx51 = (1'd0 + (4 * 32'd25));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx51_reg <= main_entry_arrayidx51;
	end
end
assign main_entry_arrayidx52 = (1'd0 + (4 * 32'd25));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx52_reg <= main_entry_arrayidx52;
	end
end
assign main_entry_arrayidx53 = (1'd0 + (4 * 32'd26));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx53_reg <= main_entry_arrayidx53;
	end
end
assign main_entry_arrayidx54 = (1'd0 + (4 * 32'd26));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx54_reg <= main_entry_arrayidx54;
	end
end
assign main_entry_arrayidx55 = (1'd0 + (4 * 32'd27));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx55_reg <= main_entry_arrayidx55;
	end
end
assign main_entry_arrayidx56 = (1'd0 + (4 * 32'd27));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx56_reg <= main_entry_arrayidx56;
	end
end
assign main_entry_arrayidx57 = (1'd0 + (4 * 32'd28));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx57_reg <= main_entry_arrayidx57;
	end
end
assign main_entry_arrayidx58 = (1'd0 + (4 * 32'd28));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx58_reg <= main_entry_arrayidx58;
	end
end
assign main_entry_arrayidx59 = (1'd0 + (4 * 32'd29));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx59_reg <= main_entry_arrayidx59;
	end
end
assign main_entry_arrayidx60 = (1'd0 + (4 * 32'd29));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx60_reg <= main_entry_arrayidx60;
	end
end
assign main_entry_arrayidx61 = (1'd0 + (4 * 32'd30));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx61_reg <= main_entry_arrayidx61;
	end
end
assign main_entry_arrayidx62 = (1'd0 + (4 * 32'd30));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx62_reg <= main_entry_arrayidx62;
	end
end
assign main_entry_arrayidx63 = (1'd0 + (4 * 32'd31));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx63_reg <= main_entry_arrayidx63;
	end
end
assign main_entry_arrayidx64 = (1'd0 + (4 * 32'd31));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_arrayidx64_reg <= main_entry_arrayidx64;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_entry_17) & (fsm_stall == 1'd0))) begin
		main_for_cond69_preheader_j67_0342 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc76_25) & (fsm_stall == 1'd0)) & (main_for_inc76_exitcond74 == 1'd0))) */ begin
		main_for_cond69_preheader_j67_0342 = main_for_inc76_4;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_entry_17) & (fsm_stall == 1'd0))) begin
		main_for_cond69_preheader_j67_0342_reg <= main_for_cond69_preheader_j67_0342;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc76_25) & (fsm_stall == 1'd0)) & (main_for_inc76_exitcond74 == 1'd0))) begin
		main_for_cond69_preheader_j67_0342_reg <= main_for_cond69_preheader_j67_0342;
	end
end
always @(*) begin
		main_for_cond69_preheader_arrayidx72 = (1'd0 + (4 * {26'd0,main_for_cond69_preheader_j67_0342_reg}));
end
always @(*) begin
		main_for_cond69_preheader_arrayidx75 = (1'd0 + (4 * {26'd0,main_for_cond69_preheader_j67_0342_reg}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond69_preheader_18)) begin
		main_for_cond69_preheader_arrayidx75_reg <= main_for_cond69_preheader_arrayidx75;
	end
end
always @(*) begin
		main_for_cond69_preheader_0 = main_entry_vla319_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond69_preheader_19)) begin
		main_for_cond69_preheader_0_reg <= main_for_cond69_preheader_0;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond69_preheader_19) & (fsm_stall == 1'd0))) begin
		main_for_body71_1 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_24) & (fsm_stall == 1'd0)) & (main_for_inc_exitcond72 == 1'd0))) */ begin
		main_for_body71_1 = main_for_inc_3;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond69_preheader_19) & (fsm_stall == 1'd0))) begin
		main_for_body71_1_reg <= main_for_body71_1;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_24) & (fsm_stall == 1'd0)) & (main_for_inc_exitcond72 == 1'd0))) begin
		main_for_body71_1_reg <= main_for_body71_1;
	end
end
always @(*) begin
		main_for_body71_arrayidx73 = (1'd0 + (4 * main_for_body71_1_reg));
end
always @(*) begin
		main_for_body71_2 = main_grid_out_a;
end
always @(*) begin
		main_for_body71_cmp74 = (main_for_cond69_preheader_0_reg == main_for_body71_2);
end
always @(*) begin
		main_for_inc_3 = (main_for_body71_1_reg + 32'd1);
end
always @(*) begin
		main_for_inc_exitcond72 = (main_for_inc_3 == 32'd36);
end
always @(*) begin
		main_for_inc76_4 = ({1'd0,main_for_cond69_preheader_j67_0342_reg} + 32'd1);
end
always @(*) begin
		main_for_inc76_exitcond74 = (main_for_inc76_4 == 32'd32);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond84_preheader_preheader_26) & (fsm_stall == 1'd0))) begin
		main_for_cond84_preheader_j79_0340 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc96_34) & (fsm_stall == 1'd0)) & (main_for_inc96_exitcond69 == 1'd0))) */ begin
		main_for_cond84_preheader_j79_0340 = main_for_inc96_9;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond84_preheader_preheader_26) & (fsm_stall == 1'd0))) begin
		main_for_cond84_preheader_j79_0340_reg <= main_for_cond84_preheader_j79_0340;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc96_34) & (fsm_stall == 1'd0)) & (main_for_inc96_exitcond69 == 1'd0))) begin
		main_for_cond84_preheader_j79_0340_reg <= main_for_cond84_preheader_j79_0340;
	end
end
always @(*) begin
		main_for_cond84_preheader_arrayidx87 = (1'd0 + (4 * {26'd0,main_for_cond84_preheader_j79_0340_reg}));
end
always @(*) begin
		main_for_cond84_preheader_arrayidx91 = (1'd0 + (4 * {26'd0,main_for_cond84_preheader_j79_0340_reg}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond84_preheader_27)) begin
		main_for_cond84_preheader_arrayidx91_reg <= main_for_cond84_preheader_arrayidx91;
	end
end
always @(*) begin
		main_for_cond84_preheader_5 = main_entry_vla1320_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond84_preheader_28)) begin
		main_for_cond84_preheader_5_reg <= main_for_cond84_preheader_5;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond84_preheader_28) & (fsm_stall == 1'd0))) begin
		main_for_body86_6 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc93_33) & (fsm_stall == 1'd0)) & (main_for_inc93_exitcond67 == 1'd0))) */ begin
		main_for_body86_6 = main_for_inc93_8;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond84_preheader_28) & (fsm_stall == 1'd0))) begin
		main_for_body86_6_reg <= main_for_body86_6;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc93_33) & (fsm_stall == 1'd0)) & (main_for_inc93_exitcond67 == 1'd0))) begin
		main_for_body86_6_reg <= main_for_body86_6;
	end
end
always @(*) begin
		main_for_body86_arrayidx88 = (1'd0 + (4 * main_for_body86_6_reg));
end
always @(*) begin
		main_for_body86_7 = main_grid_out_a;
end
always @(*) begin
		main_for_body86_cmp89 = (main_for_cond84_preheader_5_reg == main_for_body86_7);
end
always @(*) begin
		main_for_inc93_8 = (main_for_body86_6_reg + 32'd1);
end
always @(*) begin
		main_for_inc93_exitcond67 = (main_for_inc93_8 == 32'd36);
end
always @(*) begin
		main_for_inc96_9 = ({1'd0,main_for_cond84_preheader_j79_0340_reg} + 32'd1);
end
always @(*) begin
		main_for_inc96_exitcond69 = (main_for_inc96_9 == 32'd32);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body101_preheader_35) & (fsm_stall == 1'd0))) begin
		main_for_body101_i_0338 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc112_41) & (fsm_stall == 1'd0)) & (main_for_inc112_exitcond63 == 1'd0))) */ begin
		main_for_body101_i_0338 = main_for_inc112_12;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body101_preheader_35) & (fsm_stall == 1'd0))) begin
		main_for_body101_i_0338_reg <= main_for_body101_i_0338;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc112_41) & (fsm_stall == 1'd0)) & (main_for_inc112_exitcond63 == 1'd0))) begin
		main_for_body101_i_0338_reg <= main_for_body101_i_0338;
	end
end
always @(*) begin
		main_for_body101_bit_select15 = main_for_body101_i_0338_reg_width_extended[29:0];
end
always @(*) begin
		main_for_body101_bit_select13 = main_for_body101_i_0338_reg_width_extended[26:0];
end
always @(*) begin
		main_for_body101_bit_concat16 = {main_for_body101_bit_select15[29:0], main_for_body101_bit_concat16_bit_select_operand_2[1:0]};
end
always @(*) begin
		main_for_body101_bit_concat14 = {main_for_body101_bit_select13[26:0], main_for_body101_bit_concat14_bit_select_operand_2[4:0]};
end
always @(*) begin
		main_for_body101_sr_add = (main_for_body101_bit_concat16 + main_for_body101_bit_concat14);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body101_36)) begin
		main_for_body101_sr_add_reg <= main_for_body101_sr_add;
	end
end
always @(*) begin
		main_for_body101_arrayidx102 = (1'd0 + (4 * {26'd0,main_for_body101_i_0338_reg}));
end
always @(*) begin
		main_for_body101_arrayidx103 = (1'd0 + (4 * {26'd0,main_for_body101_i_0338_reg}));
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body101_37) & (fsm_stall == 1'd0))) begin
		main_for_body106_j_0337 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body106_40) & (fsm_stall == 1'd0)) & (main_for_body106_exitcond61_reg == 1'd0))) */ begin
		main_for_body106_j_0337 = main_for_body106_11_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body101_37) & (fsm_stall == 1'd0))) begin
		main_for_body106_j_0337_reg <= main_for_body106_j_0337;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body106_40) & (fsm_stall == 1'd0)) & (main_for_body106_exitcond61_reg == 1'd0))) begin
		main_for_body106_j_0337_reg <= main_for_body106_j_0337;
	end
end
always @(*) begin
		main_for_body106_10 = (main_for_body101_sr_add_reg + main_for_body106_j_0337_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body106_38)) begin
		main_for_body106_10_reg <= main_for_body106_10;
	end
end
always @(*) begin
		main_for_body106_scevgep43 = (1'd0 + (4 * main_for_body106_10_reg));
end
always @(*) begin
		main_for_body106_11 = (main_for_body106_j_0337_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body106_38)) begin
		main_for_body106_11_reg <= main_for_body106_11;
	end
end
always @(*) begin
		main_for_body106_exitcond61 = (main_for_body106_11 == 32'd36);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body106_38)) begin
		main_for_body106_exitcond61_reg <= main_for_body106_exitcond61;
	end
end
always @(*) begin
		main_for_inc112_12 = ({1'd0,main_for_body101_i_0338_reg} + 32'd1);
end
always @(*) begin
		main_for_inc112_exitcond63 = (main_for_inc112_12 == 32'd36);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond118_preheader_preheader_42) & (fsm_stall == 1'd0))) begin
		main_for_cond118_preheader_13 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc192_48) & (fsm_stall == 1'd0)) & (main_for_inc192_exitcond15 == 1'd0))) */ begin
		main_for_cond118_preheader_13 = main_for_inc192_23;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond118_preheader_preheader_42) & (fsm_stall == 1'd0))) begin
		main_for_cond118_preheader_13_reg <= main_for_cond118_preheader_13;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc192_48) & (fsm_stall == 1'd0)) & (main_for_inc192_exitcond15 == 1'd0))) begin
		main_for_cond118_preheader_13_reg <= main_for_cond118_preheader_13;
	end
end
always @(*) begin
		main_for_cond118_preheader_bit_select9 = main_for_cond118_preheader_13_reg_width_extended[26:0];
end
always @(*) begin
		main_for_cond118_preheader_bit_select7 = main_for_cond118_preheader_13_reg_width_extended[25:0];
end
always @(*) begin
		main_for_cond118_preheader_bit_select5 = main_for_cond118_preheader_13_reg_width_extended[24:0];
end
always @(*) begin
		main_for_cond118_preheader_sr_negate = (32'd0 - {1'd0,main_for_cond118_preheader_13_reg});
end
always @(*) begin
		main_for_cond118_preheader_bit_select11 = main_for_cond118_preheader_sr_negate_width_extended[30:0];
end
always @(*) begin
		main_for_cond118_preheader_bit_concat12 = {main_for_cond118_preheader_bit_select11[30:0], main_for_cond118_preheader_bit_concat12_bit_select_operand_2};
end
always @(*) begin
		main_for_cond118_preheader_bit_concat10 = {main_for_cond118_preheader_bit_select9[26:0], main_for_cond118_preheader_bit_concat10_bit_select_operand_2[4:0]};
end
always @(*) begin
		main_for_cond118_preheader_bit_concat8 = {main_for_cond118_preheader_bit_select7[25:0], main_for_cond118_preheader_bit_concat8_bit_select_operand_2[5:0]};
end
always @(*) begin
		main_for_cond118_preheader_bit_concat6 = {main_for_cond118_preheader_bit_select5[24:0], main_for_cond118_preheader_bit_concat6_bit_select_operand_2[6:0]};
end
always @(*) begin
		main_for_cond118_preheader_sr_add82 = (main_for_cond118_preheader_bit_concat12 + main_for_cond118_preheader_bit_concat10);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_43)) begin
		main_for_cond118_preheader_sr_add82_reg <= main_for_cond118_preheader_sr_add82;
	end
end
always @(*) begin
		main_for_cond118_preheader_sr_add83 = (main_for_cond118_preheader_bit_concat8 + main_for_cond118_preheader_bit_concat6);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_43)) begin
		main_for_cond118_preheader_sr_add83_reg <= main_for_cond118_preheader_sr_add83;
	end
end
always @(*) begin
		main_for_cond118_preheader_sr_add84 = (main_for_cond118_preheader_sr_add82_reg + main_for_cond118_preheader_sr_add83_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_sr_add84_reg <= main_for_cond118_preheader_sr_add84;
	end
end
always @(*) begin
		main_for_cond118_preheader_bit_select3 = main_for_cond118_preheader_sr_add84[31:1];
end
always @(*) begin
		main_for_cond118_preheader_14 = (main_for_cond118_preheader_sr_add84 + 32'd36);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_14_reg <= main_for_cond118_preheader_14;
	end
end
always @(*) begin
		main_for_cond118_preheader_scevgep41 = (1'd0 + (4 * main_for_cond118_preheader_14_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_for_cond118_preheader_scevgep41_reg <= main_for_cond118_preheader_scevgep41;
	end
end
always @(*) begin
		main_for_cond118_preheader_15 = (main_for_cond118_preheader_sr_add84 + 32'd73);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_15_reg <= main_for_cond118_preheader_15;
	end
end
always @(*) begin
		main_for_cond118_preheader_scevgep39 = (1'd0 + (4 * main_for_cond118_preheader_15_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_for_cond118_preheader_scevgep39_reg <= main_for_cond118_preheader_scevgep39;
	end
end
always @(*) begin
		main_for_cond118_preheader_16 = (main_for_cond118_preheader_sr_add84 + 32'd149);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_16_reg <= main_for_cond118_preheader_16;
	end
end
always @(*) begin
		main_for_cond118_preheader_scevgep37 = (1'd0 + (4 * main_for_cond118_preheader_16_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_for_cond118_preheader_scevgep37_reg <= main_for_cond118_preheader_scevgep37;
	end
end
always @(*) begin
		main_for_cond118_preheader_17 = (main_for_cond118_preheader_sr_add84 + 32'd184);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_17_reg <= main_for_cond118_preheader_17;
	end
end
always @(*) begin
		main_for_cond118_preheader_scevgep36 = (1'd0 + (4 * main_for_cond118_preheader_17_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_for_cond118_preheader_scevgep36_reg <= main_for_cond118_preheader_scevgep36;
	end
end
always @(*) begin
		main_for_cond118_preheader_18 = (main_for_cond118_preheader_sr_add84 + 32'd112);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_18_reg <= main_for_cond118_preheader_18;
	end
end
always @(*) begin
		main_for_cond118_preheader_scevgep35 = (1'd0 + (4 * main_for_cond118_preheader_18_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_for_cond118_preheader_scevgep35_reg <= main_for_cond118_preheader_scevgep35;
	end
end
always @(*) begin
		main_for_cond118_preheader_19 = (main_for_cond118_preheader_sr_add84 + 32'd147);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_19_reg <= main_for_cond118_preheader_19;
	end
end
always @(*) begin
		main_for_cond118_preheader_scevgep34 = (1'd0 + (4 * main_for_cond118_preheader_19_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_for_cond118_preheader_scevgep34_reg <= main_for_cond118_preheader_scevgep34;
	end
end
always @(*) begin
		main_for_cond118_preheader_20 = (main_for_cond118_preheader_sr_add84 + 32'd75);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_20_reg <= main_for_cond118_preheader_20;
	end
end
always @(*) begin
		main_for_cond118_preheader_scevgep33 = (1'd0 + (4 * main_for_cond118_preheader_20_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_for_cond118_preheader_scevgep33_reg <= main_for_cond118_preheader_scevgep33;
	end
end
always @(*) begin
		main_for_cond118_preheader_21 = (main_for_cond118_preheader_sr_add84 + 32'd110);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_21_reg <= main_for_cond118_preheader_21;
	end
end
always @(*) begin
		main_for_cond118_preheader_scevgep32 = (1'd0 + (4 * main_for_cond118_preheader_21_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_for_cond118_preheader_scevgep32_reg <= main_for_cond118_preheader_scevgep32;
	end
end
always @(*) begin
		main_for_cond118_preheader_22 = (main_for_cond118_preheader_sr_add84 + 32'd38);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_22_reg <= main_for_cond118_preheader_22;
	end
end
always @(*) begin
		main_for_cond118_preheader_scevgep31 = (1'd0 + (4 * main_for_cond118_preheader_22_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_for_cond118_preheader_scevgep31_reg <= main_for_cond118_preheader_scevgep31;
	end
end
always @(*) begin
		main_for_cond118_preheader_bit_concat4 = {main_for_cond118_preheader_bit_select3[30:0], main_for_cond118_preheader_bit_concat4_bit_select_operand_2};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_44)) begin
		main_for_cond118_preheader_bit_concat4_reg <= main_for_cond118_preheader_bit_concat4;
	end
end
always @(*) begin
		main_for_cond118_preheader_scevgep40 = (1'd0 + (4 * main_for_cond118_preheader_bit_concat4_reg));
end
always @(*) begin
		main_for_cond118_preheader_cmp121 = ($signed({28'd0,main_for_cond118_preheader_cmp121_op0_temp}) < $signed({27'd0,main_for_cond118_preheader_cmp121_op1_temp}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_43)) begin
		main_for_cond118_preheader_cmp121_reg <= main_for_cond118_preheader_cmp121;
	end
end
always @(*) begin
		main_for_inc192_23 = ({1'd0,main_for_cond118_preheader_13_reg} + 32'd1);
end
always @(*) begin
		main_for_inc192_exitcond15 = (main_for_inc192_23 == 32'd6);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body198_preheader_49) & (fsm_stall == 1'd0))) begin
		main_for_body198_i_2333 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc238_83) & (fsm_stall == 1'd0)) & (main_for_inc238_cmp196 == 1'd1))) */ begin
		main_for_body198_i_2333 = main_for_body198_inc239_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body198_preheader_49) & (fsm_stall == 1'd0))) begin
		main_for_body198_i_2333_reg <= main_for_body198_i_2333;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc238_83) & (fsm_stall == 1'd0)) & (main_for_inc238_cmp196 == 1'd1))) begin
		main_for_body198_i_2333_reg <= main_for_body198_i_2333;
	end
end
always @(*) begin
		main_for_body198_arrayidx199 = (1'd0 + (4 * {26'd0,main_for_body198_i_2333_reg}));
end
always @(*) begin
		main_for_body198_arrayidx200 = (1'd0 + (4 * {26'd0,main_for_body198_i_2333_reg}));
end
always @(*) begin
		main_for_body198_inc239 = ({1'd0,main_for_body198_i_2333_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body198_50)) begin
		main_for_body198_inc239_reg <= main_for_body198_inc239;
	end
end
always @(*) begin
		main_for_body198_24 = main_entry_vla65321_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body198_51)) begin
		main_for_body198_24_reg <= main_for_body198_24;
	end
end
always @(*) begin
		main_for_body198_25 = main_entry_vla66322_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body198_51)) begin
		main_for_body198_25_reg <= main_for_body198_25;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body198_51) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_057_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_body_i_53) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond2_reg == 1'd0))) */ begin
		main_for_body_i_i_057_i = main_for_body_i_26_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body198_51) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_057_i_reg <= main_for_body_i_i_057_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_53) & (fsm_stall == 1'd0)) & (main_for_body_i_exitcond2_reg == 1'd0))) begin
		main_for_body_i_i_057_i_reg <= main_for_body_i_i_057_i;
	end
end
always @(*) begin
		main_for_body_i_arrayidx1_i = (1'd0 + (4 * main_for_body_i_i_057_i_reg));
end
always @(*) begin
		main_for_body_i_arrayidx2_i = (1'd0 + (4 * main_for_body_i_i_057_i_reg));
end
always @(*) begin
		main_for_body_i_26 = (main_for_body_i_i_057_i_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_52)) begin
		main_for_body_i_26_reg <= main_for_body_i_26;
	end
end
always @(*) begin
		main_for_body_i_exitcond2 = (main_for_body_i_26 == 32'd36);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body_i_52)) begin
		main_for_body_i_exitcond2_reg <= main_for_body_i_exitcond2;
	end
end
always @(*) begin
		main_for_end_i_arrayidx_i = (1'd0 + (4 * main_for_body198_24_reg));
end
always @(*) begin
		main_for_end_i_arrayidx3_i = (1'd0 + (4 * main_for_body198_24_reg));
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_end_i_55) & (fsm_stall == 1'd0))) begin
		main_for_body6_i_count_056_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc31_i_74) & (fsm_stall == 1'd0)) & (main_for_inc31_i_exitcond == 1'd0))) */ begin
		main_for_body6_i_count_056_i = main_for_inc31_i_37;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_end_i_55) & (fsm_stall == 1'd0))) begin
		main_for_body6_i_count_056_i_reg <= main_for_body6_i_count_056_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc31_i_74) & (fsm_stall == 1'd0)) & (main_for_inc31_i_exitcond == 1'd0))) begin
		main_for_body6_i_count_056_i_reg <= main_for_body6_i_count_056_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_56) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_27 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_61) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond5 == 1'd0))) */ begin
		main_for_body_i_i_27 = main_for_inc_i_i_30;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_56) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_27_reg <= main_for_body_i_i_27;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_61) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond5 == 1'd0))) begin
		main_for_body_i_i_27_reg <= main_for_body_i_i_27;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_56) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_index_012_i_i = 0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_61) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond5 == 1'd0))) */ begin
		main_for_body_i_i_min_index_012_i_i = main_for_inc_i_i_min_index_1_i_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_56) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_index_012_i_i_reg <= main_for_body_i_i_min_index_012_i_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_61) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond5 == 1'd0))) begin
		main_for_body_i_i_min_index_012_i_i_reg <= main_for_body_i_i_min_index_012_i_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_56) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_011_i_i = 32'd2147483647;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_61) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond5 == 1'd0))) */ begin
		main_for_body_i_i_min_011_i_i = main_for_inc_i_i_min_1_i_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_56) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_011_i_i_reg <= main_for_body_i_i_min_011_i_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_61) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond5 == 1'd0))) begin
		main_for_body_i_i_min_011_i_i_reg <= main_for_body_i_i_min_011_i_i;
	end
end
always @(*) begin
		main_for_body_i_i_arrayidx_i_i = (1'd0 + (4 * main_for_body_i_i_27_reg));
end
always @(*) begin
		main_for_body_i_i_28 = main_entry_sptSet_i_out_a;
end
always @(*) begin
		main_for_body_i_i_cmp1_i_i = (main_for_body_i_i_28 == 32'd0);
end
always @(*) begin
		main_land_lhs_true_i_i_arrayidx2_i_i = (1'd0 + (4 * main_for_body_i_i_27_reg));
end
always @(*) begin
		main_land_lhs_true_i_i_29 = main_entry_dist_i_out_a;
end
always @(*) begin
		main_land_lhs_true_i_i_cmp3_i_i = ($signed(main_land_lhs_true_i_i_29) > $signed(main_for_body_i_i_min_011_i_i_reg));
end
always @(*) begin
		main_land_lhs_true_i_i_min_0_i_i = (main_land_lhs_true_i_i_cmp3_i_i ? main_for_body_i_i_min_011_i_i_reg : main_land_lhs_true_i_i_29);
end
always @(*) begin
		main_land_lhs_true_i_i_min_index_0_v_0_i_i = (main_land_lhs_true_i_i_cmp3_i_i ? main_for_body_i_i_min_index_012_i_i_reg : main_for_body_i_i_27_reg);
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_58) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_1_i_i = main_for_body_i_i_min_011_i_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_60) & (fsm_stall == 1'd0))) */ begin
		main_for_inc_i_i_min_1_i_i = main_land_lhs_true_i_i_min_0_i_i;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_58) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_1_i_i_reg <= main_for_inc_i_i_min_1_i_i;
	end
	if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_60) & (fsm_stall == 1'd0))) begin
		main_for_inc_i_i_min_1_i_i_reg <= main_for_inc_i_i_min_1_i_i;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_58) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_index_1_i_i = main_for_body_i_i_min_index_012_i_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_60) & (fsm_stall == 1'd0))) */ begin
		main_for_inc_i_i_min_index_1_i_i = main_land_lhs_true_i_i_min_index_0_v_0_i_i;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_58) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_index_1_i_i_reg <= main_for_inc_i_i_min_index_1_i_i;
	end
	if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_60) & (fsm_stall == 1'd0))) begin
		main_for_inc_i_i_min_index_1_i_i_reg <= main_for_inc_i_i_min_index_1_i_i;
	end
end
always @(*) begin
		main_for_inc_i_i_bit_select1 = main_for_inc_i_i_min_index_1_i_i_reg[29:0];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc_i_i_61)) begin
		main_for_inc_i_i_bit_select1_reg <= main_for_inc_i_i_bit_select1;
	end
end
always @(*) begin
		main_for_inc_i_i_bit_select = main_for_inc_i_i_min_index_1_i_i_reg[26:0];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc_i_i_61)) begin
		main_for_inc_i_i_bit_select_reg <= main_for_inc_i_i_bit_select;
	end
end
always @(*) begin
		main_for_inc_i_i_30 = (main_for_body_i_i_27_reg + 32'd1);
end
always @(*) begin
		main_for_inc_i_i_exitcond5 = (main_for_inc_i_i_30 == 32'd36);
end
always @(*) begin
		main_minDistance_exit_i_arrayidx8_i = (1'd0 + (4 * main_for_inc_i_i_min_index_1_i_i_reg));
end
always @(*) begin
		main_minDistance_exit_i_arrayidx17_i = (1'd0 + (4 * main_for_inc_i_i_min_index_1_i_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_62)) begin
		main_minDistance_exit_i_arrayidx17_i_reg <= main_minDistance_exit_i_arrayidx17_i;
	end
end
always @(*) begin
		main_minDistance_exit_i_bit_concat2 = {main_for_inc_i_i_bit_select1_reg[29:0], main_minDistance_exit_i_bit_concat2_bit_select_operand_2[1:0]};
end
always @(*) begin
		main_minDistance_exit_i_bit_concat = {main_for_inc_i_i_bit_select_reg[26:0], main_minDistance_exit_i_bit_concat_bit_select_operand_2[4:0]};
end
always @(*) begin
		main_minDistance_exit_i_sr_add87 = (main_minDistance_exit_i_bit_concat2 + main_minDistance_exit_i_bit_concat);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_62)) begin
		main_minDistance_exit_i_sr_add87_reg <= main_minDistance_exit_i_sr_add87;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_minDistance_exit_i_63) & (fsm_stall == 1'd0))) begin
		main_for_body11_i_v_055_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc28_i_73) & (fsm_stall == 1'd0)) & (main_for_inc28_i_exitcond8 == 1'd0))) */ begin
		main_for_body11_i_v_055_i = main_for_inc28_i_36;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_minDistance_exit_i_63) & (fsm_stall == 1'd0))) begin
		main_for_body11_i_v_055_i_reg <= main_for_body11_i_v_055_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc28_i_73) & (fsm_stall == 1'd0)) & (main_for_inc28_i_exitcond8 == 1'd0))) begin
		main_for_body11_i_v_055_i_reg <= main_for_body11_i_v_055_i;
	end
end
always @(*) begin
		main_for_body11_i_arrayidx12_i = (1'd0 + (4 * main_for_body11_i_v_055_i_reg));
end
always @(*) begin
		main_for_body11_i_arrayidx20_i = (1'd0 + (4 * main_for_body11_i_v_055_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body11_i_64)) begin
		main_for_body11_i_arrayidx20_i_reg <= main_for_body11_i_arrayidx20_i;
	end
end
always @(*) begin
		main_for_body11_i_arrayidx22_i = (1'd0 + (4 * main_for_body11_i_v_055_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body11_i_64)) begin
		main_for_body11_i_arrayidx22_i_reg <= main_for_body11_i_arrayidx22_i;
	end
end
always @(*) begin
		main_for_body11_i_31 = main_entry_sptSet_i_out_a;
end
always @(*) begin
		main_for_body11_i_tobool_i = (main_for_body11_i_31 == 32'd0);
end
always @(*) begin
		main_land_lhs_true_i_32 = (main_minDistance_exit_i_sr_add87_reg + main_for_body11_i_v_055_i_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_66)) begin
		main_land_lhs_true_i_32_reg <= main_land_lhs_true_i_32;
	end
end
always @(*) begin
		main_land_lhs_true_i_scevgep = (1'd0 + (4 * main_land_lhs_true_i_32_reg));
end
always @(*) begin
		main_land_lhs_true_i_33 = main_entry_m1_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_68)) begin
		main_land_lhs_true_i_33_reg <= main_land_lhs_true_i_33;
	end
end
always @(*) begin
		main_land_lhs_true_i_tobool15_i = (main_land_lhs_true_i_33 == 32'd0);
end
always @(*) begin
		main_land_lhs_true16_i_34 = main_entry_dist_i_out_a;
end
always @(*) begin
		main_land_lhs_true16_i_add_i = (main_land_lhs_true16_i_34 + main_land_lhs_true_i_33_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true16_i_70)) begin
		main_land_lhs_true16_i_add_i_reg <= main_land_lhs_true16_i_add_i;
	end
end
always @(*) begin
		main_land_lhs_true16_i_35 = main_entry_dist_i_out_b;
end
always @(*) begin
		main_land_lhs_true16_i_cmp21_i = ($signed(main_land_lhs_true16_i_add_i) < $signed(main_land_lhs_true16_i_35));
end
always @(*) begin
		main_for_inc28_i_36 = (main_for_body11_i_v_055_i_reg + 32'd1);
end
always @(*) begin
		main_for_inc28_i_exitcond8 = (main_for_inc28_i_36 == 32'd36);
end
always @(*) begin
		main_for_inc31_i_37 = (main_for_body6_i_count_056_i_reg + 32'd1);
end
always @(*) begin
		main_for_inc31_i_exitcond = (main_for_inc31_i_37 == 32'd35);
end
always @(*) begin
		main_dijkstra_exit_arrayidx207329 = (1'd0 + (4 * main_for_body198_25_reg));
end
always @(*) begin
		main_dijkstra_exit_38 = main_entry_parent_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_dijkstra_exit_76)) begin
		main_dijkstra_exit_38_reg <= main_dijkstra_exit_38;
	end
end
always @(*) begin
		main_dijkstra_exit_cmp208330 = (main_dijkstra_exit_38 == $signed(-32'd1));
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_end211_preheader_77) & (fsm_stall == 1'd0))) begin
		main_if_end211_39 = main_dijkstra_exit_38_reg;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_if_then220_81) & (fsm_stall == 1'd0)) & (main_if_then220_cmp208 == 1'd0))) */ begin
		main_if_end211_39 = main_if_then220_42;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_end211_preheader_77) & (fsm_stall == 1'd0))) begin
		main_if_end211_39_reg <= main_if_end211_39;
	end
	if ((((cur_state == LEGUP_F_main_BB_if_then220_81) & (fsm_stall == 1'd0)) & (main_if_then220_cmp208 == 1'd0))) begin
		main_if_end211_39_reg <= main_if_end211_39;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_end211_preheader_77) & (fsm_stall == 1'd0))) begin
		main_if_end211_origem_1332 = main_for_body198_25_reg;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_if_then220_81) & (fsm_stall == 1'd0)) & (main_if_then220_cmp208 == 1'd0))) */ begin
		main_if_end211_origem_1332 = main_if_end211_39_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_end211_preheader_77) & (fsm_stall == 1'd0))) begin
		main_if_end211_origem_1332_reg <= main_if_end211_origem_1332;
	end
	if ((((cur_state == LEGUP_F_main_BB_if_then220_81) & (fsm_stall == 1'd0)) & (main_if_then220_cmp208 == 1'd0))) begin
		main_if_end211_origem_1332_reg <= main_if_end211_origem_1332;
	end
end
always @(*) begin
		main_if_end211_arrayidx212 = (1'd0 + (4 * main_if_end211_39_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end211_78)) begin
		main_if_end211_arrayidx212_reg <= main_if_end211_arrayidx212;
	end
end
always @(*) begin
		main_if_end211_40 = main_entry_indice_s_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end211_79)) begin
		main_if_end211_40_reg <= main_if_end211_40;
	end
end
always @(*) begin
		main_if_end211_cmp213 = ($signed(main_if_end211_40) < $signed({27'd0,main_if_end211_cmp213_op1_temp}));
end
always @(*) begin
		main_if_end211_arrayidx215 = (1'd0 + (4 * main_if_end211_origem_1332_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end211_78)) begin
		main_if_end211_arrayidx215_reg <= main_if_end211_arrayidx215;
	end
end
always @(*) begin
		main_if_end211_41 = main_entry_indice_e_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end211_79)) begin
		main_if_end211_41_reg <= main_if_end211_41;
	end
end
always @(*) begin
		main_if_end211_cmp216 = ($signed(main_if_end211_41) < $signed({27'd0,main_if_end211_cmp216_op1_temp}));
end
always @(*) begin
		main_if_end211_and218323 = (main_if_end211_cmp213 & main_if_end211_cmp216);
end
always @(*) begin
		main_if_then220_add228 = (main_if_end211_41_reg + 32'd1);
end
always @(*) begin
		main_if_then220_add230 = (main_if_end211_40_reg + 32'd1);
end
always @(*) begin
		main_if_then220_arrayidx207 = (1'd0 + (4 * main_if_end211_39_reg));
end
always @(*) begin
		main_if_then220_42 = main_entry_parent_out_a;
end
always @(*) begin
		main_if_then220_cmp208 = (main_if_then220_42 == $signed(-32'd1));
end
always @(*) begin
		main_for_inc238_cmp196 = ($signed({24'd0,main_for_inc238_cmp196_op0_temp}) < $signed({24'd0,main_for_inc238_cmp196_op1_temp}));
end
always @(*) begin
		main_for_inc189_us_5_43 = (main_for_cond118_preheader_sr_add84_reg + 32'd253);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_43_reg <= main_for_inc189_us_5_43;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep38 = (1'd0 + (4 * main_for_inc189_us_5_43_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep38_reg <= main_for_inc189_us_5_scevgep38;
	end
end
always @(*) begin
		main_for_inc189_us_5_44 = (main_for_cond118_preheader_sr_add84_reg + 32'd401);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_44_reg <= main_for_inc189_us_5_44;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep30 = (1'd0 + (4 * main_for_inc189_us_5_44_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep30_reg <= main_for_inc189_us_5_scevgep30;
	end
end
always @(*) begin
		main_for_inc189_us_5_45 = (main_for_cond118_preheader_sr_add84_reg + 32'd191);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_45_reg <= main_for_inc189_us_5_45;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep29 = (1'd0 + (4 * main_for_inc189_us_5_45_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep29_reg <= main_for_inc189_us_5_scevgep29;
	end
end
always @(*) begin
		main_for_inc189_us_5_46 = (main_for_cond118_preheader_sr_add84_reg + 32'd364);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_46_reg <= main_for_inc189_us_5_46;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep28 = (1'd0 + (4 * main_for_inc189_us_5_46_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep28_reg <= main_for_inc189_us_5_scevgep28;
	end
end
always @(*) begin
		main_for_inc189_us_5_47 = (main_for_cond118_preheader_sr_add84_reg + 32'd154);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_47_reg <= main_for_inc189_us_5_47;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep27 = (1'd0 + (4 * main_for_inc189_us_5_47_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep27_reg <= main_for_inc189_us_5_scevgep27;
	end
end
always @(*) begin
		main_for_inc189_us_5_48 = (main_for_cond118_preheader_sr_add84_reg + 32'd327);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_48_reg <= main_for_inc189_us_5_48;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep26 = (1'd0 + (4 * main_for_inc189_us_5_48_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep26_reg <= main_for_inc189_us_5_scevgep26;
	end
end
always @(*) begin
		main_for_inc189_us_5_49 = (main_for_cond118_preheader_sr_add84_reg + 32'd117);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_49_reg <= main_for_inc189_us_5_49;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep25 = (1'd0 + (4 * main_for_inc189_us_5_49_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep25_reg <= main_for_inc189_us_5_scevgep25;
	end
end
always @(*) begin
		main_for_inc189_us_5_50 = (main_for_cond118_preheader_sr_add84_reg + 32'd290);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_50_reg <= main_for_inc189_us_5_50;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep24 = (1'd0 + (4 * main_for_inc189_us_5_50_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep24_reg <= main_for_inc189_us_5_scevgep24;
	end
end
always @(*) begin
		main_for_inc189_us_5_51 = (main_for_cond118_preheader_sr_add84_reg + 32'd80);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_51_reg <= main_for_inc189_us_5_51;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep23 = (1'd0 + (4 * main_for_inc189_us_5_51_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep23_reg <= main_for_inc189_us_5_scevgep23;
	end
end
always @(*) begin
		main_for_inc189_us_5_52 = (main_for_cond118_preheader_sr_add84_reg + 32'd43);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_52_reg <= main_for_inc189_us_5_52;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep22 = (1'd0 + (4 * main_for_inc189_us_5_52_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep22_reg <= main_for_inc189_us_5_scevgep22;
	end
end
always @(*) begin
		main_for_inc189_us_5_53 = (main_for_cond118_preheader_sr_add84_reg + 32'd216);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_53_reg <= main_for_inc189_us_5_53;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep21 = (1'd0 + (4 * main_for_inc189_us_5_53_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep21_reg <= main_for_inc189_us_5_scevgep21;
	end
end
always @(*) begin
		main_for_inc189_us_5_54 = (main_for_cond118_preheader_sr_add84_reg + 32'd6);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_for_inc189_us_5_54_reg <= main_for_inc189_us_5_54;
	end
end
always @(*) begin
		main_for_inc189_us_5_scevgep20 = (1'd0 + (4 * main_for_inc189_us_5_54_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_for_inc189_us_5_scevgep20_reg <= main_for_inc189_us_5_scevgep20;
	end
end
always @(*) begin
	main_grid_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body71_20)) begin
		main_grid_address_a = (main_for_body71_arrayidx73 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body86_29)) begin
		main_grid_address_a = (main_for_body86_arrayidx88 >>> 3'd2);
	end
end
assign main_grid_address_b = 'dx;
always @(*) begin
	main_entry_dist_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_52)) begin
		main_entry_dist_i_address_a = (main_for_body_i_arrayidx1_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_end_i_54)) begin
		main_entry_dist_i_address_a = (main_for_end_i_arrayidx3_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_59)) begin
		main_entry_dist_i_address_a = (main_land_lhs_true_i_i_arrayidx2_i_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true16_i_69)) begin
		main_entry_dist_i_address_a = (main_minDistance_exit_i_arrayidx17_i_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_dist_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_52)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end_i_54)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_dist_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_52)) begin
		main_entry_dist_i_in_a = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end_i_54)) begin
		main_entry_dist_i_in_a = 32'd0;
	end
end
always @(*) begin
	main_entry_dist_i_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true16_i_69)) begin
		main_entry_dist_i_address_b = (main_for_body11_i_arrayidx20_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_71)) begin
		main_entry_dist_i_address_b = (main_for_body11_i_arrayidx20_i_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_dist_i_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_if_then_i_71)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_dist_i_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then_i_71)) begin
		main_entry_dist_i_in_b = main_land_lhs_true16_i_add_i_reg;
	end
end
always @(*) begin
	main_entry_sptSet_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_52)) begin
		main_entry_sptSet_i_address_a = (main_for_body_i_arrayidx2_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_i_57)) begin
		main_entry_sptSet_i_address_a = (main_for_body_i_i_arrayidx_i_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_62)) begin
		main_entry_sptSet_i_address_a = (main_minDistance_exit_i_arrayidx8_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body11_i_64)) begin
		main_entry_sptSet_i_address_a = (main_for_body11_i_arrayidx12_i >>> 3'd2);
	end
end
always @(*) begin
	main_entry_sptSet_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_52)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_62)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_sptSet_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body_i_52)) begin
		main_entry_sptSet_i_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_62)) begin
		main_entry_sptSet_i_in_a = 32'd1;
	end
end
always @(*) begin
	main_entry_parent_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_end_i_54)) begin
		main_entry_parent_address_a = (main_for_end_i_arrayidx_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_71)) begin
		main_entry_parent_address_a = (main_for_body11_i_arrayidx22_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_dijkstra_exit_75)) begin
		main_entry_parent_address_a = (main_dijkstra_exit_arrayidx207329 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then220_80)) begin
		main_entry_parent_address_a = (main_if_then220_arrayidx207 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_parent_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_end_i_54)) begin
		main_entry_parent_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_71)) begin
		main_entry_parent_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_parent_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_end_i_54)) begin
		main_entry_parent_in_a = -32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_71)) begin
		main_entry_parent_in_a = main_for_inc_i_i_min_index_1_i_i_reg;
	end
end
always @(*) begin
	main_entry_m1_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body106_39)) begin
		main_entry_m1_address_a = (main_for_body106_scevgep43 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_entry_m1_address_a = (main_for_cond118_preheader_scevgep40 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_46)) begin
		main_entry_m1_address_a = (main_for_cond118_preheader_scevgep41_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_67)) begin
		main_entry_m1_address_a = (main_land_lhs_true_i_scevgep >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_87)) begin
		main_entry_m1_address_a = (main_for_cond118_preheader_scevgep31_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_88)) begin
		main_entry_m1_address_a = (main_for_cond118_preheader_scevgep33_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_89)) begin
		main_entry_m1_address_a = (main_for_cond118_preheader_scevgep35_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_90)) begin
		main_entry_m1_address_a = (main_for_cond118_preheader_scevgep37_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_entry_m1_address_a = (main_for_cond118_preheader_scevgep31_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_entry_m1_address_a = (main_for_cond118_preheader_scevgep33_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_94)) begin
		main_entry_m1_address_a = (main_for_cond118_preheader_scevgep35_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_95)) begin
		main_entry_m1_address_a = (main_for_cond118_preheader_scevgep37_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_96)) begin
		main_entry_m1_address_a = (main_for_inc189_us_5_scevgep20_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_97)) begin
		main_entry_m1_address_a = (main_for_inc189_us_5_scevgep22_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_98)) begin
		main_entry_m1_address_a = (main_for_inc189_us_5_scevgep23_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_99)) begin
		main_entry_m1_address_a = (main_for_inc189_us_5_scevgep25_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_100)) begin
		main_entry_m1_address_a = (main_for_inc189_us_5_scevgep27_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_101)) begin
		main_entry_m1_address_a = (main_for_inc189_us_5_scevgep29_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_m1_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body106_39)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_46)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_87)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_88)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_89)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_90)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_94)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_95)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_96)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_97)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_98)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_99)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_100)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_101)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_m1_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body106_39)) begin
		main_entry_m1_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_45)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond118_preheader_46)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_87)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_88)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_89)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_90)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_94)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_95)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_96)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_97)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_98)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_99)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_100)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_101)) begin
		main_entry_m1_in_a = 32'd1;
	end
end
always @(*) begin
	main_entry_m1_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_87)) begin
		main_entry_m1_address_b = (main_for_cond118_preheader_scevgep39_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_88)) begin
		main_entry_m1_address_b = (main_for_cond118_preheader_scevgep32_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_89)) begin
		main_entry_m1_address_b = (main_for_cond118_preheader_scevgep34_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_90)) begin
		main_entry_m1_address_b = (main_for_cond118_preheader_scevgep36_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_entry_m1_address_b = (main_for_cond118_preheader_scevgep39_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_entry_m1_address_b = (main_for_cond118_preheader_scevgep32_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_94)) begin
		main_entry_m1_address_b = (main_for_cond118_preheader_scevgep34_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_95)) begin
		main_entry_m1_address_b = (main_for_cond118_preheader_scevgep36_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_96)) begin
		main_entry_m1_address_b = (main_for_inc189_us_5_scevgep21_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_97)) begin
		main_entry_m1_address_b = (main_for_inc189_us_5_scevgep38_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_98)) begin
		main_entry_m1_address_b = (main_for_inc189_us_5_scevgep24_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_99)) begin
		main_entry_m1_address_b = (main_for_inc189_us_5_scevgep26_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_100)) begin
		main_entry_m1_address_b = (main_for_inc189_us_5_scevgep28_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_101)) begin
		main_entry_m1_address_b = (main_for_inc189_us_5_scevgep30_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_m1_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_87)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_88)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_89)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_90)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_94)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_95)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_96)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_97)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_98)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_99)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_100)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_101)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_m1_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_87)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_88)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_89)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_5_90)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_92)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_93)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_94)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_95)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_96)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_97)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_98)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_99)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_100)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc189_us_5_101)) begin
		main_entry_m1_in_b = 32'd1;
	end
end
always @(*) begin
	main_entry_indice_e_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body101_36)) begin
		main_entry_indice_e_address_a = (main_for_body101_arrayidx102 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end211_78)) begin
		main_entry_indice_e_address_a = (main_if_end211_arrayidx215 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then220_80)) begin
		main_entry_indice_e_address_a = (main_if_end211_arrayidx215_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_indice_e_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body101_36)) begin
		main_entry_indice_e_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then220_80)) begin
		main_entry_indice_e_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_indice_e_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body101_36)) begin
		main_entry_indice_e_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then220_80)) begin
		main_entry_indice_e_in_a = main_if_then220_add228;
	end
end
always @(*) begin
	main_entry_indice_s_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body101_36)) begin
		main_entry_indice_s_address_a = (main_for_body101_arrayidx103 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end211_78)) begin
		main_entry_indice_s_address_a = (main_if_end211_arrayidx212 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then220_80)) begin
		main_entry_indice_s_address_a = (main_if_end211_arrayidx212_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_indice_s_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body101_36)) begin
		main_entry_indice_s_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then220_80)) begin
		main_entry_indice_s_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_indice_s_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body101_36)) begin
		main_entry_indice_s_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then220_80)) begin
		main_entry_indice_s_in_a = main_if_then220_add230;
	end
end
always @(*) begin
	main_entry_vla319_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla319_address_a = (main_entry_vla319_sub >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx5_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx9_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx13_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx17_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx21_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx25_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx29_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx33_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx37_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx41_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx45_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx49_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx53_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx57_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla319_address_a = (main_entry_arrayidx61_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond69_preheader_18)) begin
		main_entry_vla319_address_a = (main_for_cond69_preheader_arrayidx72 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla319_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla319_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla319_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla319_in_a = 32'd26;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla319_in_a = 32'd25;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla319_in_a = 32'd23;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla319_in_a = 32'd20;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla319_in_a = 32'd15;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla319_in_a = 32'd9;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla319_in_a = 32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla319_in_a = 32'd7;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla319_in_a = 32'd11;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla319_in_a = 32'd21;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla319_in_a = 32'd17;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla319_in_a = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla319_in_a = 32'd24;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla319_in_a = 32'd19;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla319_in_a = 32'd12;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla319_in_a = 32'd14;
	end
end
always @(*) begin
	main_entry_vla319_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx3 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx7_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx11_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx15_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx19_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx23_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx27_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx31_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx35_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx39_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx43_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx47_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx51_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx55_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx59_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla319_address_b = (main_entry_arrayidx63_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla319_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla319_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_vla319_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla319_in_b = 32'd25;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla319_in_b = 32'd23;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla319_in_b = 32'd20;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla319_in_b = 32'd15;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla319_in_b = 32'd9;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla319_in_b = 32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla319_in_b = 32'd13;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla319_in_b = 32'd18;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla319_in_b = 32'd21;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla319_in_b = 32'd17;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla319_in_b = 32'd10;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla319_in_b = 32'd16;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla319_in_b = 32'd22;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla319_in_b = 32'd19;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla319_in_b = 32'd6;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla319_in_b = 32'd8;
	end
end
always @(*) begin
	main_entry_vla1320_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1320_address_a = (main_entry_vla1320_sub >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx6_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx10_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx14_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx18_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx22_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx26_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx30_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx34_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx38_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx42_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx46_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx50_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx54_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx58_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1320_address_a = (main_entry_arrayidx62_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond84_preheader_27)) begin
		main_entry_vla1320_address_a = (main_for_cond84_preheader_arrayidx87 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla1320_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1320_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla1320_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1320_in_a = 32'd25;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1320_in_a = 32'd23;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1320_in_a = 32'd20;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1320_in_a = 32'd15;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1320_in_a = 32'd9;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1320_in_a = 32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1320_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1320_in_a = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1320_in_a = 32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1320_in_a = 32'd17;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1320_in_a = 32'd13;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1320_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1320_in_a = 32'd22;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1320_in_a = 32'd14;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1320_in_a = 32'd6;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1320_in_a = 32'd8;
	end
end
always @(*) begin
	main_entry_vla1320_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx4 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx8_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx12_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx16_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx20_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx24_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx28_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx32_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx36_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx40_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx44_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx48_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx52_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx56_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx60_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1320_address_b = (main_entry_arrayidx64_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla1320_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1320_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_vla1320_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla1320_in_b = 32'd24;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla1320_in_b = 32'd21;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla1320_in_b = 32'd18;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla1320_in_b = 32'd13;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla1320_in_b = 32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla1320_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla1320_in_b = 32'd7;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla1320_in_b = 32'd11;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla1320_in_b = 32'd16;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_10)) begin
		main_entry_vla1320_in_b = 32'd10;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_11)) begin
		main_entry_vla1320_in_b = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_12)) begin
		main_entry_vla1320_in_b = 32'd10;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_13)) begin
		main_entry_vla1320_in_b = 32'd19;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_14)) begin
		main_entry_vla1320_in_b = 32'd12;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_15)) begin
		main_entry_vla1320_in_b = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_16)) begin
		main_entry_vla1320_in_b = 32'd2;
	end
end
always @(*) begin
	main_entry_vla65321_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then_22)) begin
		main_entry_vla65321_address_a = (main_for_cond69_preheader_arrayidx75_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body198_50)) begin
		main_entry_vla65321_address_a = (main_for_body198_arrayidx199 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla65321_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_if_then_22)) begin
		main_entry_vla65321_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla65321_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then_22)) begin
		main_entry_vla65321_in_a = main_for_body71_1_reg;
	end
end
always @(*) begin
	main_entry_vla66322_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then90_31)) begin
		main_entry_vla66322_address_a = (main_for_cond84_preheader_arrayidx91_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body198_50)) begin
		main_entry_vla66322_address_a = (main_for_body198_arrayidx200 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla66322_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_if_then90_31)) begin
		main_entry_vla66322_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla66322_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_if_then90_31)) begin
		main_entry_vla66322_in_a = main_for_body86_6_reg;
	end
end
always @(*) begin
	main_for_body101_i_0338_reg_width_extended = {24'd0,main_for_body101_i_0338_reg};
end
assign main_for_body101_bit_concat16_bit_select_operand_2 = 2'd0;
assign main_for_body101_bit_concat14_bit_select_operand_2 = 5'd0;
always @(*) begin
	main_for_cond118_preheader_13_reg_width_extended = {24'd0,main_for_cond118_preheader_13_reg};
end
always @(*) begin
	main_for_cond118_preheader_sr_negate_width_extended = {{27{main_for_cond118_preheader_sr_negate[3]}},main_for_cond118_preheader_sr_negate};
end
assign main_for_cond118_preheader_bit_concat12_bit_select_operand_2 = 1'd0;
assign main_for_cond118_preheader_bit_concat10_bit_select_operand_2 = 5'd0;
assign main_for_cond118_preheader_bit_concat8_bit_select_operand_2 = 6'd0;
assign main_for_cond118_preheader_bit_concat6_bit_select_operand_2 = 7'd0;
always @(*) begin
	main_for_cond118_preheader_cmp121_op0_temp = {1'd0,main_for_cond118_preheader_13_reg};
end
assign main_for_cond118_preheader_cmp121_op1_temp = 32'd5;
assign main_for_cond118_preheader_bit_concat4_bit_select_operand_2 = 1'd1;
assign main_minDistance_exit_i_bit_concat2_bit_select_operand_2 = 2'd0;
assign main_minDistance_exit_i_bit_concat_bit_select_operand_2 = 5'd0;
assign main_if_end211_cmp213_op1_temp = 32'd4;
assign main_if_end211_cmp216_op1_temp = 32'd4;
always @(*) begin
	main_for_inc238_cmp196_op0_temp = {1'd0,main_for_body198_inc239_reg};
end
assign main_for_inc238_cmp196_op1_temp = 32'd32;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end240_86)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end240_86)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "Arria10",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module ram_single_port_intel
(
	clk,
	clken,
	address_a,
	wren_a,
	data_a,
	byteena_a,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
    .wren_a (wren_a),
    .data_a (data_a),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.operation_mode = "SINGLE_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "Arria10",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module rom_dual_port
(
	clk,
	clken,
	address_a,
	q_a,
	address_b,
	q_b
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  init_file = {`MEM_INIT_DIR, "UNUSED.mif"};
parameter  latency = 1;

input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
reg [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
reg [(width_b-1):0] q_b_wire;

(* ram_init_file = init_file *) reg [width_a-1:0] ram [numwords_a-1:0];

integer i;
/* synthesis translate_off */
ALTERA_MF_MEMORY_INITIALIZATION mem ();
reg [8*256:1] ram_ver_file;
initial begin
	if (init_file == {`MEM_INIT_DIR, "UNUSED.mif"})
    begin
		for (i = 0; i < numwords_a; i = i + 1)
			ram[i] = 0;
    end
	else
    begin
        // modelsim can't read .mif files directly. So use Altera function to
        // convert them to .ver files
        mem.convert_to_ver_file(init_file, width_a, ram_ver_file);
        $readmemh(ram_ver_file, ram);
    end
end
/* synthesis translate_on */

localparam input_latency = ((latency - 1) >> 1);
localparam output_latency = (latency - 1) - input_latency;
integer j;

reg [(widthad_a-1):0] address_a_reg[input_latency:0];
reg [(widthad_b-1):0] address_b_reg[input_latency:0];

always @(*)
begin
  address_a_reg[0] = address_a;
  address_b_reg[0] = address_b;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < input_latency; j=j+1)
   begin
       address_a_reg[j+1] <= address_a_reg[j];
       address_b_reg[j+1] <= address_b_reg[j];
   end
end

always @ (posedge clk)
if (clken)
begin
    q_a_wire <= ram[address_a_reg[input_latency]];
end

always @ (posedge clk)
if (clken)
begin
    q_b_wire <= ram[address_b_reg[input_latency]];
end


reg [(width_a-1):0] q_a_reg[output_latency:0];

always @(*)
begin
   q_a_reg[0] <= q_a_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_a_reg[j+1] <= q_a_reg[j];
   end
end

assign q_a = q_a_reg[output_latency];
reg [(width_b-1):0] q_b_reg[output_latency:0];

always @(*)
begin
   q_b_reg[0] <= q_b_wire;
end

always @(posedge clk)
if (clken)
begin
   for (j = 0; j < output_latency; j=j+1)
   begin
       q_b_reg[j+1] <= q_b_reg[j];
   end
end

assign q_b = q_b_reg[output_latency];

endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
