// ----------------------------------------------------------------------------
// LegUp High-Level Synthesis Tool Version 7.5 (http://legupcomputing.com)
// Copyright (c) 2015-2019 LegUp Computing Inc. All Rights Reserved.
// For technical issues, please contact: support@legupcomputing.com
// For general inquiries, please contact: info@legupcomputing.com
// Date: Fri May  8 21:41:58 2020
// ----------------------------------------------------------------------------
`define MEMORY_CONTROLLER_ADDR_SIZE 32
// This directory contains the memory initialization files generated by LegUp.
// This relative path is used by ModelSim and FPGA synthesis tool.
`define MEM_INIT_DIR "../mem_init/"

`timescale 1 ns / 1 ns
module top
(
	clk,
	reset,
	start,
	finish,
	return_val
);

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg  main_inst_clk;
reg  main_inst_reset;
reg  main_inst_start;
wire  main_inst_finish;
wire [31:0] main_inst_return_val;
reg  main_inst_finish_reg;
reg [31:0] main_inst_return_val_reg;


main main_inst (
	.clk (main_inst_clk),
	.reset (main_inst_reset),
	.start (main_inst_start),
	.finish (main_inst_finish),
	.return_val (main_inst_return_val)
);



always @(*) begin
	main_inst_clk = clk;
end
always @(*) begin
	main_inst_reset = reset;
end
always @(*) begin
	main_inst_start = start;
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_finish_reg <= 1'd0;
	end
	if (main_inst_finish) begin
		main_inst_finish_reg <= 1'd1;
	end
end
always @(posedge clk) begin
	if ((reset | main_inst_start)) begin
		main_inst_return_val_reg <= 0;
	end
	if (main_inst_finish) begin
		main_inst_return_val_reg <= main_inst_return_val;
	end
end
always @(*) begin
	finish = main_inst_finish;
end
always @(*) begin
	return_val = main_inst_return_val;
end

endmodule
`timescale 1 ns / 1 ns
module main
(
	clk,
	reset,
	start,
	finish,
	return_val
);

parameter [7:0] LEGUP_0 = 8'd0;
parameter [7:0] LEGUP_F_main_BB_entry_1 = 8'd1;
parameter [7:0] LEGUP_F_main_BB_entry_2 = 8'd2;
parameter [7:0] LEGUP_F_main_BB_entry_3 = 8'd3;
parameter [7:0] LEGUP_F_main_BB_entry_4 = 8'd4;
parameter [7:0] LEGUP_F_main_BB_entry_5 = 8'd5;
parameter [7:0] LEGUP_F_main_BB_entry_6 = 8'd6;
parameter [7:0] LEGUP_F_main_BB_entry_7 = 8'd7;
parameter [7:0] LEGUP_F_main_BB_entry_8 = 8'd8;
parameter [7:0] LEGUP_F_main_BB_entry_9 = 8'd9;
parameter [7:0] LEGUP_F_main_BB_entry_10 = 8'd10;
parameter [7:0] LEGUP_F_main_BB_for_cond43_preheader_11 = 8'd11;
parameter [7:0] LEGUP_F_main_BB_NodeBlock27_12 = 8'd12;
parameter [7:0] LEGUP_F_main_BB_NodeBlock25_13 = 8'd13;
parameter [7:0] LEGUP_F_main_BB_NodeBlock23_14 = 8'd14;
parameter [7:0] LEGUP_F_main_BB_LeafBlock21_15 = 8'd15;
parameter [7:0] LEGUP_F_main_BB_NodeBlock19_16 = 8'd16;
parameter [7:0] LEGUP_F_main_BB_NodeBlock17_17 = 8'd17;
parameter [7:0] LEGUP_F_main_BB_NodeBlock15_18 = 8'd18;
parameter [7:0] LEGUP_F_main_BB_NodeBlock13_19 = 8'd19;
parameter [7:0] LEGUP_F_main_BB_NodeBlock11_20 = 8'd20;
parameter [7:0] LEGUP_F_main_BB_NodeBlock9_21 = 8'd21;
parameter [7:0] LEGUP_F_main_BB_NodeBlock7_22 = 8'd22;
parameter [7:0] LEGUP_F_main_BB_NodeBlock5_23 = 8'd23;
parameter [7:0] LEGUP_F_main_BB_NodeBlock3_24 = 8'd24;
parameter [7:0] LEGUP_F_main_BB_NodeBlock1_25 = 8'd25;
parameter [7:0] LEGUP_F_main_BB_NodeBlock_26 = 8'd26;
parameter [7:0] LEGUP_F_main_BB_LeafBlock_27 = 8'd27;
parameter [7:0] LEGUP_F_main_BB_for_cond58_preheader_28 = 8'd28;
parameter [7:0] LEGUP_F_main_BB_NodeBlock62_29 = 8'd29;
parameter [7:0] LEGUP_F_main_BB_NodeBlock60_30 = 8'd30;
parameter [7:0] LEGUP_F_main_BB_NodeBlock58_31 = 8'd31;
parameter [7:0] LEGUP_F_main_BB_LeafBlock56_32 = 8'd32;
parameter [7:0] LEGUP_F_main_BB_NodeBlock54_33 = 8'd33;
parameter [7:0] LEGUP_F_main_BB_NodeBlock52_34 = 8'd34;
parameter [7:0] LEGUP_F_main_BB_NodeBlock50_35 = 8'd35;
parameter [7:0] LEGUP_F_main_BB_NodeBlock48_36 = 8'd36;
parameter [7:0] LEGUP_F_main_BB_NodeBlock46_37 = 8'd37;
parameter [7:0] LEGUP_F_main_BB_NodeBlock44_38 = 8'd38;
parameter [7:0] LEGUP_F_main_BB_NodeBlock42_39 = 8'd39;
parameter [7:0] LEGUP_F_main_BB_NodeBlock40_40 = 8'd40;
parameter [7:0] LEGUP_F_main_BB_NodeBlock38_41 = 8'd41;
parameter [7:0] LEGUP_F_main_BB_NodeBlock36_42 = 8'd42;
parameter [7:0] LEGUP_F_main_BB_NodeBlock34_43 = 8'd43;
parameter [7:0] LEGUP_F_main_BB_LeafBlock32_44 = 8'd44;
parameter [7:0] LEGUP_F_main_BB_for_body75_45 = 8'd45;
parameter [7:0] LEGUP_F_main_BB_for_body75_46 = 8'd46;
parameter [7:0] LEGUP_F_main_BB_for_body75_47 = 8'd47;
parameter [7:0] LEGUP_F_main_BB_for_body75_48 = 8'd48;
parameter [7:0] LEGUP_F_main_BB_for_body75_49 = 8'd49;
parameter [7:0] LEGUP_F_main_BB_for_body75_50 = 8'd50;
parameter [7:0] LEGUP_F_main_BB_for_body75_51 = 8'd51;
parameter [7:0] LEGUP_F_main_BB_for_body75_52 = 8'd52;
parameter [7:0] LEGUP_F_main_BB_for_body75_53 = 8'd53;
parameter [7:0] LEGUP_F_main_BB_for_body75_54 = 8'd54;
parameter [7:0] LEGUP_F_main_BB_for_body75_55 = 8'd55;
parameter [7:0] LEGUP_F_main_BB_for_body75_56 = 8'd56;
parameter [7:0] LEGUP_F_main_BB_for_body75_57 = 8'd57;
parameter [7:0] LEGUP_F_main_BB_for_body75_58 = 8'd58;
parameter [7:0] LEGUP_F_main_BB_for_body75_59 = 8'd59;
parameter [7:0] LEGUP_F_main_BB_for_body75_60 = 8'd60;
parameter [7:0] LEGUP_F_main_BB_for_body75_61 = 8'd61;
parameter [7:0] LEGUP_F_main_BB_for_cond92_preheader_preheader_62 = 8'd62;
parameter [7:0] LEGUP_F_main_BB_for_cond92_preheader_63 = 8'd63;
parameter [7:0] LEGUP_F_main_BB_for_cond92_preheader_64 = 8'd64;
parameter [7:0] LEGUP_F_main_BB_for_cond92_preheader_65 = 8'd65;
parameter [7:0] LEGUP_F_main_BB_for_cond92_preheader_66 = 8'd66;
parameter [7:0] LEGUP_F_main_BB_for_cond169_preheader_67 = 8'd67;
parameter [7:0] LEGUP_F_main_BB_for_inc166_68 = 8'd68;
parameter [7:0] LEGUP_F_main_BB_for_body172_69 = 8'd69;
parameter [7:0] LEGUP_F_main_BB_for_body172_70 = 8'd70;
parameter [7:0] LEGUP_F_main_BB_for_body172_71 = 8'd71;
parameter [7:0] LEGUP_F_main_BB_for_body172_72 = 8'd72;
parameter [7:0] LEGUP_F_main_BB_for_body172_73 = 8'd73;
parameter [7:0] LEGUP_F_main_BB_for_body172_74 = 8'd74;
parameter [7:0] LEGUP_F_main_BB_for_body172_75 = 8'd75;
parameter [7:0] LEGUP_F_main_BB_for_body172_76 = 8'd76;
parameter [7:0] LEGUP_F_main_BB_for_body172_77 = 8'd77;
parameter [7:0] LEGUP_F_main_BB_for_body172_78 = 8'd78;
parameter [7:0] LEGUP_F_main_BB_for_body6_i_79 = 8'd79;
parameter [7:0] LEGUP_F_main_BB_for_body_i_i_80 = 8'd80;
parameter [7:0] LEGUP_F_main_BB_for_body_i_i_81 = 8'd81;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true_i_i_82 = 8'd82;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true_i_i_83 = 8'd83;
parameter [7:0] LEGUP_F_main_BB_for_inc_i_i_84 = 8'd84;
parameter [7:0] LEGUP_F_main_BB_minDistance_exit_i_85 = 8'd85;
parameter [7:0] LEGUP_F_main_BB_minDistance_exit_i_86 = 8'd86;
parameter [7:0] LEGUP_F_main_BB_for_body11_i_87 = 8'd87;
parameter [7:0] LEGUP_F_main_BB_for_body11_i_88 = 8'd88;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true_i_89 = 8'd89;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true_i_90 = 8'd90;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true_i_91 = 8'd91;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true16_i_92 = 8'd92;
parameter [7:0] LEGUP_F_main_BB_land_lhs_true16_i_93 = 8'd93;
parameter [7:0] LEGUP_F_main_BB_if_then_i_94 = 8'd94;
parameter [7:0] LEGUP_F_main_BB_if_then_i_95 = 8'd95;
parameter [7:0] LEGUP_F_main_BB_for_inc28_i_96 = 8'd96;
parameter [7:0] LEGUP_F_main_BB_for_inc31_i_97 = 8'd97;
parameter [7:0] LEGUP_F_main_BB_dijkstra_exit_98 = 8'd98;
parameter [7:0] LEGUP_F_main_BB_dijkstra_exit_99 = 8'd99;
parameter [7:0] LEGUP_F_main_BB_if_end185_preheader_100 = 8'd100;
parameter [7:0] LEGUP_F_main_BB_if_end185_101 = 8'd101;
parameter [7:0] LEGUP_F_main_BB_if_end185_102 = 8'd102;
parameter [7:0] LEGUP_F_main_BB_if_then194_103 = 8'd103;
parameter [7:0] LEGUP_F_main_BB_if_then194_104 = 8'd104;
parameter [7:0] LEGUP_F_main_BB_for_inc212_loopexit_105 = 8'd105;
parameter [7:0] LEGUP_F_main_BB_for_inc212_106 = 8'd106;
parameter [7:0] LEGUP_F_main_BB_for_end214_loopexit_107 = 8'd107;
parameter [7:0] LEGUP_F_main_BB_for_end214_loopexit1_108 = 8'd108;
parameter [7:0] LEGUP_F_main_BB_for_end214_109 = 8'd109;
parameter [7:0] LEGUP_F_main_BB_for_inc163_3_110 = 8'd110;
parameter [7:0] LEGUP_F_main_BB_for_inc163_3_111 = 8'd111;
parameter [7:0] LEGUP_F_main_BB_for_inc163_3_112 = 8'd112;
parameter [7:0] LEGUP_F_main_BB_for_inc163_us_3_113 = 8'd113;
parameter [7:0] LEGUP_F_main_BB_for_inc163_us_3_114 = 8'd114;
parameter [7:0] LEGUP_F_main_BB_for_inc163_us_3_115 = 8'd115;
parameter [7:0] LEGUP_F_main_BB_for_inc163_us_3_116 = 8'd116;
parameter [7:0] LEGUP_F_main_BB_for_inc163_us_3_117 = 8'd117;
parameter [7:0] LEGUP_F_main_BB_for_inc163_us_3_118 = 8'd118;
parameter [7:0] LEGUP_F_main_BB_for_inc163_us_3_119 = 8'd119;
parameter [7:0] LEGUP_F_main_BB_for_inc67_15_storemerge_120 = 8'd120;
parameter [7:0] LEGUP_F_main_BB_for_inc67_15_storemerge_121 = 8'd121;
parameter [7:0] LEGUP_F_main_BB_for_inc67_15_122 = 8'd122;
parameter [7:0] LEGUP_F_main_BB_for_body75_preheader_123 = 8'd123;
parameter [7:0] LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_124 = 8'd124;
parameter [7:0] LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_125 = 8'd125;
parameter [7:0] LEGUP_F_main_BB_for_inc_15_storemerge_126 = 8'd126;
parameter [7:0] LEGUP_F_main_BB_for_inc_15_storemerge_127 = 8'd127;
parameter [7:0] LEGUP_F_main_BB_for_inc_15_128 = 8'd128;
parameter [7:0] LEGUP_F_main_BB_for_cond58_preheader_preheader_129 = 8'd129;
parameter [7:0] LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_130 = 8'd130;
parameter [7:0] LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_131 = 8'd131;

input  clk;
input  reset;
input  start;
output reg  finish;
output reg [31:0] return_val;
reg [7:0] cur_state/* synthesis syn_encoding="onehot" */;
reg [7:0] next_state;
wire  fsm_stall;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_0;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_1;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_2;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_3;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_4;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_4_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_5;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_5_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_6;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_6_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_7;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_7_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_8;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_8_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_9;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_9_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_10;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_10_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_11;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_11_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_12;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_12_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_13;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_13_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_14;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_14_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_15;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_15_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_16;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_16_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_17;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_17_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_18;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_18_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_19;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_19_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_20;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_20_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_21;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_21_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_22;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_22_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_23;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_23_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_24;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_24_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_25;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_25_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_26;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_26_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_27;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_27_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_28;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_28_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_29;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_29_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_30;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_30_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_31;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_31_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_32;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_32_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_33;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_33_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_34;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_34_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_35;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_entry_35_reg;
reg [31:0] main_for_cond43_preheader_36;
reg [31:0] main_for_cond43_preheader_36_reg;
reg [31:0] main_for_cond43_preheader_37;
reg [31:0] main_for_cond43_preheader_37_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond43_preheader_arrayidx49;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond43_preheader_arrayidx49_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond43_preheader_scevgep49;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond43_preheader_scevgep49_reg;
reg [31:0] main_for_cond43_preheader_38;
reg [31:0] main_for_cond43_preheader_38_reg;
reg  main_for_cond43_preheader_Pivot30;
reg  main_NodeBlock27_Pivot28;
reg  main_NodeBlock25_Pivot26;
reg  main_NodeBlock23_Pivot24;
reg  main_LeafBlock21_SwitchLeaf22;
reg  main_NodeBlock19_Pivot20;
reg [3:0] main_NodeBlock19_1;
reg  main_NodeBlock17_Pivot18;
reg  main_NodeBlock15_Pivot16;
reg [3:0] main_NodeBlock15_66;
reg  main_NodeBlock13_Pivot14;
reg [3:0] main_NodeBlock13_67;
reg  main_NodeBlock11_Pivot12;
reg  main_NodeBlock9_Pivot10;
reg  main_NodeBlock7_Pivot8;
reg [2:0] main_NodeBlock7_68;
reg  main_NodeBlock5_Pivot6;
reg [3:0] main_NodeBlock5_69;
reg  main_NodeBlock3_Pivot4;
reg  main_NodeBlock1_Pivot2;
reg [3:0] main_NodeBlock1_70;
reg  main_NodeBlock_Pivot;
reg  main_LeafBlock_SwitchLeaf;
reg [31:0] main_for_cond58_preheader_39;
reg [31:0] main_for_cond58_preheader_39_reg;
reg [31:0] main_for_cond58_preheader_40;
reg [31:0] main_for_cond58_preheader_40_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond58_preheader_arrayidx65;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond58_preheader_arrayidx65_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond58_preheader_scevgep47;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond58_preheader_scevgep47_reg;
reg [31:0] main_for_cond58_preheader_41;
reg [31:0] main_for_cond58_preheader_41_reg;
reg  main_for_cond58_preheader_Pivot65;
reg  main_NodeBlock62_Pivot63;
reg  main_NodeBlock60_Pivot61;
reg  main_NodeBlock58_Pivot59;
reg  main_LeafBlock56_SwitchLeaf57;
reg  main_NodeBlock54_Pivot55;
reg [3:0] main_NodeBlock54_71;
reg  main_NodeBlock52_Pivot53;
reg  main_NodeBlock50_Pivot51;
reg [3:0] main_NodeBlock50_72;
reg  main_NodeBlock48_Pivot49;
reg [3:0] main_NodeBlock48_73;
reg  main_NodeBlock46_Pivot47;
reg  main_NodeBlock44_Pivot45;
reg  main_NodeBlock42_Pivot43;
reg [2:0] main_NodeBlock42_74;
reg  main_NodeBlock40_Pivot41;
reg [3:0] main_NodeBlock40_75;
reg  main_NodeBlock38_Pivot39;
reg  main_NodeBlock36_Pivot37;
reg [3:0] main_NodeBlock36_76;
reg  main_NodeBlock34_Pivot35;
reg  main_LeafBlock32_SwitchLeaf33;
reg [4:0] main_for_body75_i_0312;
reg [4:0] main_for_body75_i_0312_reg;
reg [27:0] main_for_body75_bit_select7;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_arrayidx76;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_arrayidx77;
reg [31:0] main_for_body75_bit_concat23;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep44;
reg [31:0] main_for_body75_bit_concat22;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep43;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep43_reg;
reg [31:0] main_for_body75_bit_concat21;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep42;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep42_reg;
reg [31:0] main_for_body75_bit_concat20;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep41;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep41_reg;
reg [31:0] main_for_body75_bit_concat19;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep40;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep40_reg;
reg [31:0] main_for_body75_bit_concat18;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep39;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep39_reg;
reg [31:0] main_for_body75_bit_concat17;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep38;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep38_reg;
reg [31:0] main_for_body75_bit_concat16;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep37;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep37_reg;
reg [31:0] main_for_body75_bit_concat15;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep36;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep36_reg;
reg [31:0] main_for_body75_bit_concat14;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep35;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep35_reg;
reg [31:0] main_for_body75_bit_concat13;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep34;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep34_reg;
reg [31:0] main_for_body75_bit_concat12;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep33;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep33_reg;
reg [31:0] main_for_body75_bit_concat11;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep32;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep32_reg;
reg [31:0] main_for_body75_bit_concat10;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep31;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep31_reg;
reg [31:0] main_for_body75_bit_concat9;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep30;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep30_reg;
reg [31:0] main_for_body75_bit_concat8;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep29;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body75_scevgep29_reg;
reg [5:0] main_for_body75_42;
reg [5:0] main_for_body75_42_reg;
reg  main_for_body75_exitcond59;
reg  main_for_body75_exitcond59_reg;
reg [2:0] main_for_cond92_preheader_43;
reg [2:0] main_for_cond92_preheader_43_reg;
reg [29:0] main_for_cond92_preheader_bit_select5;
reg [25:0] main_for_cond92_preheader_bit_select3;
reg [31:0] main_for_cond92_preheader_bit_concat6;
reg [31:0] main_for_cond92_preheader_bit_concat4;
reg [31:0] main_for_cond92_preheader_sr_add;
reg [31:0] main_for_cond92_preheader_sr_add_reg;
reg [30:0] main_for_cond92_preheader_bit_select1;
reg [31:0] main_for_cond92_preheader_44;
reg [31:0] main_for_cond92_preheader_44_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep27;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep27_reg;
reg [31:0] main_for_cond92_preheader_bit_concat2;
reg [31:0] main_for_cond92_preheader_bit_concat2_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep26;
reg [31:0] main_for_cond92_preheader_45;
reg [31:0] main_for_cond92_preheader_45_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep25;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep25_reg;
reg [31:0] main_for_cond92_preheader_46;
reg [31:0] main_for_cond92_preheader_46_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep23;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep23_reg;
reg [31:0] main_for_cond92_preheader_47;
reg [31:0] main_for_cond92_preheader_47_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep22;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep22_reg;
reg [31:0] main_for_cond92_preheader_48;
reg [31:0] main_for_cond92_preheader_48_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep20;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond92_preheader_scevgep20_reg;
reg  main_for_cond92_preheader_cmp95;
reg  main_for_cond92_preheader_cmp95_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_1_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_1_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_1_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_1_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_2_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_2_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_2_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_2_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_3_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_3_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_3_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_3_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_4_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_4_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_4_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_4_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_5_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_5_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_5_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_5_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_6_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_6_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_6_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_6_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_7_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_7_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_7_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_7_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_8_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_8_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_8_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_8_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_9_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_9_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_9_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_9_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_10_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_10_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_10_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_10_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_11_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_11_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_11_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_11_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_12_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_12_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_12_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_12_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_13_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_13_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_13_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_13_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_14_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_14_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_14_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_14_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_15_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx1_15_i_reg;
wire [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_15_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_cond169_preheader_arrayidx2_15_i_reg;
reg [3:0] main_for_inc166_49;
reg  main_for_inc166_exitcond12;
reg [4:0] main_for_body172_i_2307;
reg [4:0] main_for_body172_i_2307_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body172_arrayidx173;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body172_arrayidx174;
reg [5:0] main_for_body172_inc213;
reg [5:0] main_for_body172_inc213_reg;
reg [31:0] main_for_body172_50;
reg [31:0] main_for_body172_51;
reg [31:0] main_for_body172_51_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body172_arrayidx_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body172_arrayidx3_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body172_arrayidx3_i_reg;
reg [31:0] main_for_body6_i_count_056_i;
reg [31:0] main_for_body6_i_count_056_i_reg;
reg [31:0] main_for_body_i_i_52;
reg [31:0] main_for_body_i_i_52_reg;
reg [31:0] main_for_body_i_i_min_index_012_i_i;
reg [31:0] main_for_body_i_i_min_index_012_i_i_reg;
reg [31:0] main_for_body_i_i_min_011_i_i;
reg [31:0] main_for_body_i_i_min_011_i_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body_i_i_arrayidx_i_i;
reg [31:0] main_for_body_i_i_53;
reg  main_for_body_i_i_cmp1_i_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_land_lhs_true_i_i_arrayidx2_i_i;
reg [31:0] main_land_lhs_true_i_i_54;
reg  main_land_lhs_true_i_i_cmp3_i_i;
reg [31:0] main_land_lhs_true_i_i_min_0_i_i;
reg [31:0] main_land_lhs_true_i_i_min_index_0_v_0_i_i;
reg [31:0] main_for_inc_i_i_min_1_i_i;
reg [31:0] main_for_inc_i_i_min_1_i_i_reg;
reg [31:0] main_for_inc_i_i_min_index_1_i_i;
reg [31:0] main_for_inc_i_i_min_index_1_i_i_reg;
reg [27:0] main_for_inc_i_i_bit_select;
reg [27:0] main_for_inc_i_i_bit_select_reg;
reg [31:0] main_for_inc_i_i_55;
reg  main_for_inc_i_i_exitcond2;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_minDistance_exit_i_arrayidx8_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_minDistance_exit_i_arrayidx17_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_minDistance_exit_i_arrayidx17_i_reg;
reg [31:0] main_minDistance_exit_i_bit_concat;
reg [31:0] main_minDistance_exit_i_bit_concat_reg;
reg [31:0] main_for_body11_i_v_055_i;
reg [31:0] main_for_body11_i_v_055_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx12_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx20_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx20_i_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx22_i;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_body11_i_arrayidx22_i_reg;
reg [31:0] main_for_body11_i_56;
reg  main_for_body11_i_tobool_i;
reg [31:0] main_land_lhs_true_i_57;
reg [31:0] main_land_lhs_true_i_57_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_land_lhs_true_i_scevgep;
reg [31:0] main_land_lhs_true_i_58;
reg [31:0] main_land_lhs_true_i_58_reg;
reg  main_land_lhs_true_i_tobool15_i;
reg [31:0] main_land_lhs_true16_i_59;
reg [31:0] main_land_lhs_true16_i_add_i;
reg [31:0] main_land_lhs_true16_i_add_i_reg;
reg [31:0] main_land_lhs_true16_i_60;
reg  main_land_lhs_true16_i_cmp21_i;
reg [31:0] main_for_inc28_i_61;
reg  main_for_inc28_i_exitcond;
reg [31:0] main_for_inc31_i_62;
reg  main_for_inc31_i_exitcond9;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_dijkstra_exit_arrayidx181303;
reg [31:0] main_dijkstra_exit_63;
reg [31:0] main_dijkstra_exit_63_reg;
reg  main_dijkstra_exit_cmp182304;
reg [31:0] main_if_end185_64;
reg [31:0] main_if_end185_64_reg;
reg [31:0] main_if_end185_origem_1306;
reg [31:0] main_if_end185_origem_1306_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end185_arrayidx186;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end185_arrayidx186_reg;
reg [31:0] main_if_end185_65;
reg [31:0] main_if_end185_65_reg;
reg  main_if_end185_cmp187;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end185_arrayidx189;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_end185_arrayidx189_reg;
reg [31:0] main_if_end185_66;
reg [31:0] main_if_end185_66_reg;
reg  main_if_end185_cmp190;
reg  main_if_end185_and192297;
reg [31:0] main_if_then194_add202;
reg [31:0] main_if_then194_add204;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_if_then194_arrayidx181;
reg [31:0] main_if_then194_67;
reg  main_if_then194_cmp182;
reg  main_for_inc212_cmp170;
reg [31:0] main_for_inc163_us_3_68;
reg [31:0] main_for_inc163_us_3_68_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep24;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep24_reg;
reg [31:0] main_for_inc163_us_3_69;
reg [31:0] main_for_inc163_us_3_69_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep21;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep21_reg;
reg [31:0] main_for_inc163_us_3_70;
reg [31:0] main_for_inc163_us_3_70_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep19;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep19_reg;
reg [31:0] main_for_inc163_us_3_71;
reg [31:0] main_for_inc163_us_3_71_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep18;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep18_reg;
reg [31:0] main_for_inc163_us_3_72;
reg [31:0] main_for_inc163_us_3_72_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep17;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep17_reg;
reg [31:0] main_for_inc163_us_3_73;
reg [31:0] main_for_inc163_us_3_73_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep16;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep16_reg;
reg [31:0] main_for_inc163_us_3_74;
reg [31:0] main_for_inc163_us_3_74_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep15;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep15_reg;
reg [31:0] main_for_inc163_us_3_75;
reg [31:0] main_for_inc163_us_3_75_reg;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep14;
reg [`MEMORY_CONTROLLER_ADDR_SIZE-1:0] main_for_inc163_us_3_scevgep14_reg;
reg [3:0] main_for_inc67_15_storemerge_storemerge52;
reg [3:0] main_for_inc67_15_storemerge_storemerge52_reg;
reg  main_for_inc67_15_exitcond322;
reg [31:0] main_for_inc67_15_for_cond58_preheader_crit_edge_p;
reg [3:0] main_for_inc_15_storemerge_storemerge;
reg [3:0] main_for_inc_15_storemerge_storemerge_reg;
reg  main_for_inc_15_exitcond324;
reg [31:0] main_for_inc_15_for_cond43_preheader_crit_edge_pre;
reg [3:0] main_entry_dist_i_address_a;
reg  main_entry_dist_i_write_enable_a;
reg [31:0] main_entry_dist_i_in_a;
wire [31:0] main_entry_dist_i_out_a;
reg [3:0] main_entry_dist_i_address_b;
reg  main_entry_dist_i_write_enable_b;
reg [31:0] main_entry_dist_i_in_b;
wire [31:0] main_entry_dist_i_out_b;
reg [3:0] main_entry_sptSet_i_address_a;
reg  main_entry_sptSet_i_write_enable_a;
reg [31:0] main_entry_sptSet_i_in_a;
wire [31:0] main_entry_sptSet_i_out_a;
reg [3:0] main_entry_sptSet_i_address_b;
reg  main_entry_sptSet_i_write_enable_b;
reg [31:0] main_entry_sptSet_i_in_b;
wire [31:0] main_entry_sptSet_i_out_b;
reg [3:0] main_entry_parent_address_a;
reg  main_entry_parent_write_enable_a;
reg [31:0] main_entry_parent_in_a;
wire [31:0] main_entry_parent_out_a;
reg [7:0] main_entry_m1_address_a;
reg  main_entry_m1_write_enable_a;
reg [31:0] main_entry_m1_in_a;
wire [31:0] main_entry_m1_out_a;
reg [7:0] main_entry_m1_address_b;
reg  main_entry_m1_write_enable_b;
reg [31:0] main_entry_m1_in_b;
wire [31:0] main_entry_m1_out_b;
reg [3:0] main_entry_indice_e_address_a;
reg  main_entry_indice_e_write_enable_a;
reg [31:0] main_entry_indice_e_in_a;
wire [31:0] main_entry_indice_e_out_a;
reg [3:0] main_entry_indice_s_address_a;
reg  main_entry_indice_s_write_enable_a;
reg [31:0] main_entry_indice_s_in_a;
wire [31:0] main_entry_indice_s_out_a;
reg [4:0] main_entry_vla2932_address_a;
reg  main_entry_vla2932_write_enable_a;
reg [31:0] main_entry_vla2932_in_a;
wire [31:0] main_entry_vla2932_out_a;
reg [4:0] main_entry_vla2932_address_b;
reg  main_entry_vla2932_write_enable_b;
reg [31:0] main_entry_vla2932_in_b;
wire [31:0] main_entry_vla2932_out_b;
reg [4:0] main_entry_vla12943_address_a;
reg  main_entry_vla12943_write_enable_a;
reg [31:0] main_entry_vla12943_in_a;
wire [31:0] main_entry_vla12943_out_a;
reg [4:0] main_entry_vla12943_address_b;
reg  main_entry_vla12943_write_enable_b;
reg [31:0] main_entry_vla12943_in_b;
wire [31:0] main_entry_vla12943_out_b;
reg [4:0] main_entry_vla39295_address_a;
reg  main_entry_vla39295_write_enable_a;
reg [31:0] main_entry_vla39295_in_a;
wire [31:0] main_entry_vla39295_out_a;
reg [4:0] main_entry_vla40296_address_a;
reg  main_entry_vla40296_write_enable_a;
reg [31:0] main_entry_vla40296_in_a;
wire [31:0] main_entry_vla40296_out_a;
wire [5:0] main_for_cond43_preheader_Pivot30_op1_temp;
wire [5:0] main_NodeBlock27_Pivot28_op1_temp;
wire [5:0] main_NodeBlock25_Pivot26_op1_temp;
wire [5:0] main_NodeBlock23_Pivot24_op1_temp;
wire [5:0] main_NodeBlock19_Pivot20_op1_temp;
wire [5:0] main_NodeBlock17_Pivot18_op1_temp;
wire [5:0] main_NodeBlock15_Pivot16_op1_temp;
wire [5:0] main_NodeBlock13_Pivot14_op1_temp;
wire [4:0] main_NodeBlock11_Pivot12_op1_temp;
wire [4:0] main_NodeBlock9_Pivot10_op1_temp;
wire [4:0] main_NodeBlock7_Pivot8_op1_temp;
wire [4:0] main_NodeBlock5_Pivot6_op1_temp;
wire [3:0] main_NodeBlock3_Pivot4_op1_temp;
wire [3:0] main_NodeBlock1_Pivot2_op1_temp;
wire [2:0] main_NodeBlock_Pivot_op1_temp;
wire [5:0] main_for_cond58_preheader_Pivot65_op1_temp;
wire [5:0] main_NodeBlock62_Pivot63_op1_temp;
wire [5:0] main_NodeBlock60_Pivot61_op1_temp;
wire [5:0] main_NodeBlock58_Pivot59_op1_temp;
wire [5:0] main_NodeBlock54_Pivot55_op1_temp;
wire [5:0] main_NodeBlock52_Pivot53_op1_temp;
wire [5:0] main_NodeBlock50_Pivot51_op1_temp;
wire [5:0] main_NodeBlock48_Pivot49_op1_temp;
wire [4:0] main_NodeBlock46_Pivot47_op1_temp;
wire [4:0] main_NodeBlock44_Pivot45_op1_temp;
wire [4:0] main_NodeBlock42_Pivot43_op1_temp;
wire [4:0] main_NodeBlock40_Pivot41_op1_temp;
wire [3:0] main_NodeBlock38_Pivot39_op1_temp;
wire [3:0] main_NodeBlock36_Pivot37_op1_temp;
wire [2:0] main_NodeBlock34_Pivot35_op1_temp;
reg [27:0] main_for_body75_i_0312_reg_width_extended;
wire [3:0] main_for_body75_bit_concat23_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat22_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat21_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat20_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat19_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat18_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat17_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat16_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat15_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat14_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat13_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat12_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat11_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat10_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat9_bit_select_operand_2;
wire [3:0] main_for_body75_bit_concat8_bit_select_operand_2;
reg [29:0] main_for_cond92_preheader_43_reg_width_extended;
wire [1:0] main_for_cond92_preheader_bit_concat6_bit_select_operand_2;
wire [5:0] main_for_cond92_preheader_bit_concat4_bit_select_operand_2;
wire  main_for_cond92_preheader_bit_concat2_bit_select_operand_2;
reg [3:0] main_for_cond92_preheader_cmp95_op0_temp;
wire [3:0] main_for_cond92_preheader_cmp95_op1_temp;
wire [3:0] main_minDistance_exit_i_bit_concat_bit_select_operand_2;
wire [4:0] main_if_end185_cmp187_op1_temp;
wire [4:0] main_if_end185_cmp190_op1_temp;
reg [6:0] main_for_inc212_cmp170_op0_temp;
wire [6:0] main_for_inc212_cmp170_op1_temp;



//   %dist.i = alloca [16 x i32], align 4, !dbg !83, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_dist_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_dist_i_address_a ),
	.wren_a( main_entry_dist_i_write_enable_a ),
	.data_a( main_entry_dist_i_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_dist_i_out_a ),
	.address_b( main_entry_dist_i_address_b ),
	.wren_b( main_entry_dist_i_write_enable_b ),
	.data_b( main_entry_dist_i_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_dist_i_out_b )
);
defparam main_entry_dist_i.width_a = 32;
defparam main_entry_dist_i.widthad_a = 4;
defparam main_entry_dist_i.width_be_a = 4;
defparam main_entry_dist_i.numwords_a = 16;
defparam main_entry_dist_i.width_b = 32;
defparam main_entry_dist_i.widthad_b = 4;
defparam main_entry_dist_i.width_be_b = 4;
defparam main_entry_dist_i.numwords_b = 16;
defparam main_entry_dist_i.latency = 1;


//   %sptSet.i = alloca [16 x i32], align 4, !dbg !83, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_sptSet_i (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_sptSet_i_address_a ),
	.wren_a( main_entry_sptSet_i_write_enable_a ),
	.data_a( main_entry_sptSet_i_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_sptSet_i_out_a ),
	.address_b( main_entry_sptSet_i_address_b ),
	.wren_b( main_entry_sptSet_i_write_enable_b ),
	.data_b( main_entry_sptSet_i_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_sptSet_i_out_b )
);
defparam main_entry_sptSet_i.width_a = 32;
defparam main_entry_sptSet_i.widthad_a = 4;
defparam main_entry_sptSet_i.width_be_a = 4;
defparam main_entry_sptSet_i.numwords_a = 16;
defparam main_entry_sptSet_i.width_b = 32;
defparam main_entry_sptSet_i.widthad_b = 4;
defparam main_entry_sptSet_i.width_be_b = 4;
defparam main_entry_sptSet_i.numwords_b = 16;
defparam main_entry_sptSet_i.latency = 1;


//   %parent = alloca [16 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_parent (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_parent_address_a ),
	.wren_a( main_entry_parent_write_enable_a ),
	.data_a( main_entry_parent_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_parent_out_a )
);
defparam main_entry_parent.width_a = 32;
defparam main_entry_parent.widthad_a = 4;
defparam main_entry_parent.width_be_a = 4;
defparam main_entry_parent.numwords_a = 16;
defparam main_entry_parent.latency = 1;


//   %m1 = alloca [256 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_m1 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_m1_address_a ),
	.wren_a( main_entry_m1_write_enable_a ),
	.data_a( main_entry_m1_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_m1_out_a ),
	.address_b( main_entry_m1_address_b ),
	.wren_b( main_entry_m1_write_enable_b ),
	.data_b( main_entry_m1_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_m1_out_b )
);
defparam main_entry_m1.width_a = 32;
defparam main_entry_m1.widthad_a = 8;
defparam main_entry_m1.width_be_a = 4;
defparam main_entry_m1.numwords_a = 256;
defparam main_entry_m1.width_b = 32;
defparam main_entry_m1.widthad_b = 8;
defparam main_entry_m1.width_be_b = 4;
defparam main_entry_m1.numwords_b = 256;
defparam main_entry_m1.latency = 1;


//   %indice_e = alloca [16 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_indice_e (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_indice_e_address_a ),
	.wren_a( main_entry_indice_e_write_enable_a ),
	.data_a( main_entry_indice_e_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_indice_e_out_a )
);
defparam main_entry_indice_e.width_a = 32;
defparam main_entry_indice_e.widthad_a = 4;
defparam main_entry_indice_e.width_be_a = 4;
defparam main_entry_indice_e.numwords_a = 16;
defparam main_entry_indice_e.latency = 1;


//   %indice_s = alloca [16 x i32], align 4, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_indice_s (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_indice_s_address_a ),
	.wren_a( main_entry_indice_s_write_enable_a ),
	.data_a( main_entry_indice_s_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_indice_s_out_a )
);
defparam main_entry_indice_s.width_a = 32;
defparam main_entry_indice_s.widthad_a = 4;
defparam main_entry_indice_s.width_be_a = 4;
defparam main_entry_indice_s.numwords_a = 16;
defparam main_entry_indice_s.latency = 1;


//   %vla2932 = alloca [18 x i32], align 4, !dbg !88, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_vla2932 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla2932_address_a ),
	.wren_a( main_entry_vla2932_write_enable_a ),
	.data_a( main_entry_vla2932_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla2932_out_a ),
	.address_b( main_entry_vla2932_address_b ),
	.wren_b( main_entry_vla2932_write_enable_b ),
	.data_b( main_entry_vla2932_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_vla2932_out_b )
);
defparam main_entry_vla2932.width_a = 32;
defparam main_entry_vla2932.widthad_a = 5;
defparam main_entry_vla2932.width_be_a = 4;
defparam main_entry_vla2932.numwords_a = 18;
defparam main_entry_vla2932.width_b = 32;
defparam main_entry_vla2932.widthad_b = 5;
defparam main_entry_vla2932.width_be_b = 4;
defparam main_entry_vla2932.numwords_b = 18;
defparam main_entry_vla2932.latency = 1;


//   %vla12943 = alloca [18 x i32], align 4, !dbg !89, !MSB !86, !LSB !87, !extendFrom !86
ram_dual_port main_entry_vla12943 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla12943_address_a ),
	.wren_a( main_entry_vla12943_write_enable_a ),
	.data_a( main_entry_vla12943_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla12943_out_a ),
	.address_b( main_entry_vla12943_address_b ),
	.wren_b( main_entry_vla12943_write_enable_b ),
	.data_b( main_entry_vla12943_in_b ),
	.byteena_b( {4{1'b1}} ),
	.q_b( main_entry_vla12943_out_b )
);
defparam main_entry_vla12943.width_a = 32;
defparam main_entry_vla12943.widthad_a = 5;
defparam main_entry_vla12943.width_be_a = 4;
defparam main_entry_vla12943.numwords_a = 18;
defparam main_entry_vla12943.width_b = 32;
defparam main_entry_vla12943.widthad_b = 5;
defparam main_entry_vla12943.width_be_b = 4;
defparam main_entry_vla12943.numwords_b = 18;
defparam main_entry_vla12943.latency = 1;


//   %vla40296 = alloca [19 x i32], align 4, !dbg !130, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_vla40296 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla40296_address_a ),
	.wren_a( main_entry_vla40296_write_enable_a ),
	.data_a( main_entry_vla40296_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla40296_out_a )
);
defparam main_entry_vla40296.width_a = 32;
defparam main_entry_vla40296.widthad_a = 5;
defparam main_entry_vla40296.width_be_a = 4;
defparam main_entry_vla40296.numwords_a = 19;
defparam main_entry_vla40296.latency = 1;


//   %vla39295 = alloca [19 x i32], align 4, !dbg !130, !MSB !86, !LSB !87, !extendFrom !86
ram_single_port_intel main_entry_vla39295 (
	.clk( clk ),
	.clken( !fsm_stall ),
	.address_a( main_entry_vla39295_address_a ),
	.wren_a( main_entry_vla39295_write_enable_a ),
	.data_a( main_entry_vla39295_in_a ),
	.byteena_a( {4{1'b1}} ),
	.q_a( main_entry_vla39295_out_a )
);
defparam main_entry_vla39295.width_a = 32;
defparam main_entry_vla39295.widthad_a = 5;
defparam main_entry_vla39295.width_be_a = 4;
defparam main_entry_vla39295.numwords_a = 19;
defparam main_entry_vla39295.latency = 1;

always @(posedge clk) begin
if (reset == 1'b1)
	cur_state <= LEGUP_0;
else if (!fsm_stall)
	cur_state <= next_state;
end

always @(*)
begin
next_state = cur_state;
case(cur_state)  /* synthesis parallel_case */
LEGUP_0:
	if ((fsm_stall == 1'd0) && (start == 1'd1))
		next_state = LEGUP_F_main_BB_entry_1;
LEGUP_F_main_BB_LeafBlock21_15:
	if ((fsm_stall == 1'd0) && (main_LeafBlock21_SwitchLeaf22 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_126;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock21_SwitchLeaf22 == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc_15_128;
LEGUP_F_main_BB_LeafBlock32_44:
	if ((fsm_stall == 1'd0) && (main_LeafBlock32_SwitchLeaf33 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_120;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock32_SwitchLeaf33 == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc67_15_122;
LEGUP_F_main_BB_LeafBlock56_32:
	if ((fsm_stall == 1'd0) && (main_LeafBlock56_SwitchLeaf57 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_120;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock56_SwitchLeaf57 == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc67_15_122;
LEGUP_F_main_BB_LeafBlock_27:
	if ((fsm_stall == 1'd0) && (main_LeafBlock_SwitchLeaf == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_126;
	else if ((fsm_stall == 1'd0) && (main_LeafBlock_SwitchLeaf == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc_15_128;
LEGUP_F_main_BB_NodeBlock11_20:
	if ((fsm_stall == 1'd0) && (main_NodeBlock11_Pivot12 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock3_24;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock11_Pivot12 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock9_21;
LEGUP_F_main_BB_NodeBlock13_19:
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_126;
LEGUP_F_main_BB_NodeBlock15_18:
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_126;
LEGUP_F_main_BB_NodeBlock17_17:
	if ((fsm_stall == 1'd0) && (main_NodeBlock17_Pivot18 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock13_19;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock17_Pivot18 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock15_18;
LEGUP_F_main_BB_NodeBlock19_16:
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_126;
LEGUP_F_main_BB_NodeBlock1_25:
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_126;
LEGUP_F_main_BB_NodeBlock23_14:
	if ((fsm_stall == 1'd0) && (main_NodeBlock23_Pivot24 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_126;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock23_Pivot24 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock21_15;
LEGUP_F_main_BB_NodeBlock25_13:
	if ((fsm_stall == 1'd0) && (main_NodeBlock25_Pivot26 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock19_16;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock25_Pivot26 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock23_14;
LEGUP_F_main_BB_NodeBlock27_12:
	if ((fsm_stall == 1'd0) && (main_NodeBlock27_Pivot28 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock17_17;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock27_Pivot28 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock25_13;
LEGUP_F_main_BB_NodeBlock34_43:
	if ((fsm_stall == 1'd0) && (main_NodeBlock34_Pivot35 == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock32_44;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock34_Pivot35 == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_120;
LEGUP_F_main_BB_NodeBlock36_42:
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_120;
LEGUP_F_main_BB_NodeBlock38_41:
	if ((fsm_stall == 1'd0) && (main_NodeBlock38_Pivot39 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock34_43;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock38_Pivot39 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock36_42;
LEGUP_F_main_BB_NodeBlock3_24:
	if ((fsm_stall == 1'd0) && (main_NodeBlock3_Pivot4 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock_26;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock3_Pivot4 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock1_25;
LEGUP_F_main_BB_NodeBlock40_40:
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_120;
LEGUP_F_main_BB_NodeBlock42_39:
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_120;
LEGUP_F_main_BB_NodeBlock44_38:
	if ((fsm_stall == 1'd0) && (main_NodeBlock44_Pivot45 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock40_40;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock44_Pivot45 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock42_39;
LEGUP_F_main_BB_NodeBlock46_37:
	if ((fsm_stall == 1'd0) && (main_NodeBlock46_Pivot47 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock38_41;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock46_Pivot47 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock44_38;
LEGUP_F_main_BB_NodeBlock48_36:
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_120;
LEGUP_F_main_BB_NodeBlock50_35:
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_120;
LEGUP_F_main_BB_NodeBlock52_34:
	if ((fsm_stall == 1'd0) && (main_NodeBlock52_Pivot53 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock48_36;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock52_Pivot53 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock50_35;
LEGUP_F_main_BB_NodeBlock54_33:
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_120;
LEGUP_F_main_BB_NodeBlock58_31:
	if ((fsm_stall == 1'd0) && (main_NodeBlock58_Pivot59 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_120;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock58_Pivot59 == 1'd0))
		next_state = LEGUP_F_main_BB_LeafBlock56_32;
LEGUP_F_main_BB_NodeBlock5_23:
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_126;
LEGUP_F_main_BB_NodeBlock60_30:
	if ((fsm_stall == 1'd0) && (main_NodeBlock60_Pivot61 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock54_33;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock60_Pivot61 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock58_31;
LEGUP_F_main_BB_NodeBlock62_29:
	if ((fsm_stall == 1'd0) && (main_NodeBlock62_Pivot63 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock52_34;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock62_Pivot63 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock60_30;
LEGUP_F_main_BB_NodeBlock7_22:
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_126;
LEGUP_F_main_BB_NodeBlock9_21:
	if ((fsm_stall == 1'd0) && (main_NodeBlock9_Pivot10 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock5_23;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock9_Pivot10 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock7_22;
LEGUP_F_main_BB_NodeBlock_26:
	if ((fsm_stall == 1'd0) && (main_NodeBlock_Pivot == 1'd1))
		next_state = LEGUP_F_main_BB_LeafBlock_27;
	else if ((fsm_stall == 1'd0) && (main_NodeBlock_Pivot == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_126;
LEGUP_F_main_BB_dijkstra_exit_98:
		next_state = LEGUP_F_main_BB_dijkstra_exit_99;
LEGUP_F_main_BB_dijkstra_exit_99:
	if ((fsm_stall == 1'd0) && (main_dijkstra_exit_cmp182304 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc212_106;
	else if ((fsm_stall == 1'd0) && (main_dijkstra_exit_cmp182304 == 1'd0))
		next_state = LEGUP_F_main_BB_if_end185_preheader_100;
LEGUP_F_main_BB_entry_1:
		next_state = LEGUP_F_main_BB_entry_2;
LEGUP_F_main_BB_entry_10:
		next_state = LEGUP_F_main_BB_for_cond43_preheader_11;
LEGUP_F_main_BB_entry_2:
		next_state = LEGUP_F_main_BB_entry_3;
LEGUP_F_main_BB_entry_3:
		next_state = LEGUP_F_main_BB_entry_4;
LEGUP_F_main_BB_entry_4:
		next_state = LEGUP_F_main_BB_entry_5;
LEGUP_F_main_BB_entry_5:
		next_state = LEGUP_F_main_BB_entry_6;
LEGUP_F_main_BB_entry_6:
		next_state = LEGUP_F_main_BB_entry_7;
LEGUP_F_main_BB_entry_7:
		next_state = LEGUP_F_main_BB_entry_8;
LEGUP_F_main_BB_entry_8:
		next_state = LEGUP_F_main_BB_entry_9;
LEGUP_F_main_BB_entry_9:
		next_state = LEGUP_F_main_BB_entry_10;
LEGUP_F_main_BB_for_body11_i_87:
		next_state = LEGUP_F_main_BB_for_body11_i_88;
LEGUP_F_main_BB_for_body11_i_88:
	if ((fsm_stall == 1'd0) && (main_for_body11_i_tobool_i == 1'd1))
		next_state = LEGUP_F_main_BB_land_lhs_true_i_89;
	else if ((fsm_stall == 1'd0) && (main_for_body11_i_tobool_i == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc28_i_96;
LEGUP_F_main_BB_for_body172_69:
		next_state = LEGUP_F_main_BB_for_body172_70;
LEGUP_F_main_BB_for_body172_70:
		next_state = LEGUP_F_main_BB_for_body172_71;
LEGUP_F_main_BB_for_body172_71:
		next_state = LEGUP_F_main_BB_for_body172_72;
LEGUP_F_main_BB_for_body172_72:
		next_state = LEGUP_F_main_BB_for_body172_73;
LEGUP_F_main_BB_for_body172_73:
		next_state = LEGUP_F_main_BB_for_body172_74;
LEGUP_F_main_BB_for_body172_74:
		next_state = LEGUP_F_main_BB_for_body172_75;
LEGUP_F_main_BB_for_body172_75:
		next_state = LEGUP_F_main_BB_for_body172_76;
LEGUP_F_main_BB_for_body172_76:
		next_state = LEGUP_F_main_BB_for_body172_77;
LEGUP_F_main_BB_for_body172_77:
		next_state = LEGUP_F_main_BB_for_body172_78;
LEGUP_F_main_BB_for_body172_78:
		next_state = LEGUP_F_main_BB_for_body6_i_79;
LEGUP_F_main_BB_for_body6_i_79:
		next_state = LEGUP_F_main_BB_for_body_i_i_80;
LEGUP_F_main_BB_for_body75_45:
		next_state = LEGUP_F_main_BB_for_body75_46;
LEGUP_F_main_BB_for_body75_46:
		next_state = LEGUP_F_main_BB_for_body75_47;
LEGUP_F_main_BB_for_body75_47:
		next_state = LEGUP_F_main_BB_for_body75_48;
LEGUP_F_main_BB_for_body75_48:
		next_state = LEGUP_F_main_BB_for_body75_49;
LEGUP_F_main_BB_for_body75_49:
		next_state = LEGUP_F_main_BB_for_body75_50;
LEGUP_F_main_BB_for_body75_50:
		next_state = LEGUP_F_main_BB_for_body75_51;
LEGUP_F_main_BB_for_body75_51:
		next_state = LEGUP_F_main_BB_for_body75_52;
LEGUP_F_main_BB_for_body75_52:
		next_state = LEGUP_F_main_BB_for_body75_53;
LEGUP_F_main_BB_for_body75_53:
		next_state = LEGUP_F_main_BB_for_body75_54;
LEGUP_F_main_BB_for_body75_54:
		next_state = LEGUP_F_main_BB_for_body75_55;
LEGUP_F_main_BB_for_body75_55:
		next_state = LEGUP_F_main_BB_for_body75_56;
LEGUP_F_main_BB_for_body75_56:
		next_state = LEGUP_F_main_BB_for_body75_57;
LEGUP_F_main_BB_for_body75_57:
		next_state = LEGUP_F_main_BB_for_body75_58;
LEGUP_F_main_BB_for_body75_58:
		next_state = LEGUP_F_main_BB_for_body75_59;
LEGUP_F_main_BB_for_body75_59:
		next_state = LEGUP_F_main_BB_for_body75_60;
LEGUP_F_main_BB_for_body75_60:
		next_state = LEGUP_F_main_BB_for_body75_61;
LEGUP_F_main_BB_for_body75_61:
	if ((fsm_stall == 1'd0) && (main_for_body75_exitcond59_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond92_preheader_preheader_62;
	else if ((fsm_stall == 1'd0) && (main_for_body75_exitcond59_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_body75_45;
LEGUP_F_main_BB_for_body75_preheader_123:
		next_state = LEGUP_F_main_BB_for_body75_45;
LEGUP_F_main_BB_for_body_i_i_80:
		next_state = LEGUP_F_main_BB_for_body_i_i_81;
LEGUP_F_main_BB_for_body_i_i_81:
	if ((fsm_stall == 1'd0) && (main_for_body_i_i_cmp1_i_i == 1'd1))
		next_state = LEGUP_F_main_BB_land_lhs_true_i_i_82;
	else if ((fsm_stall == 1'd0) && (main_for_body_i_i_cmp1_i_i == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc_i_i_84;
LEGUP_F_main_BB_for_cond169_preheader_67:
		next_state = LEGUP_F_main_BB_for_body172_69;
LEGUP_F_main_BB_for_cond43_preheader_11:
	if ((fsm_stall == 1'd0) && (main_for_cond43_preheader_Pivot30 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock11_20;
	else if ((fsm_stall == 1'd0) && (main_for_cond43_preheader_Pivot30 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock27_12;
LEGUP_F_main_BB_for_cond58_preheader_28:
	if ((fsm_stall == 1'd0) && (main_for_cond58_preheader_Pivot65 == 1'd1))
		next_state = LEGUP_F_main_BB_NodeBlock46_37;
	else if ((fsm_stall == 1'd0) && (main_for_cond58_preheader_Pivot65 == 1'd0))
		next_state = LEGUP_F_main_BB_NodeBlock62_29;
LEGUP_F_main_BB_for_cond58_preheader_preheader_129:
		next_state = LEGUP_F_main_BB_for_cond58_preheader_28;
LEGUP_F_main_BB_for_cond92_preheader_63:
		next_state = LEGUP_F_main_BB_for_cond92_preheader_64;
LEGUP_F_main_BB_for_cond92_preheader_64:
		next_state = LEGUP_F_main_BB_for_cond92_preheader_65;
LEGUP_F_main_BB_for_cond92_preheader_65:
		next_state = LEGUP_F_main_BB_for_cond92_preheader_66;
LEGUP_F_main_BB_for_cond92_preheader_66:
	if ((fsm_stall == 1'd0) && (main_for_cond92_preheader_cmp95_reg == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc163_us_3_113;
	else if ((fsm_stall == 1'd0) && (main_for_cond92_preheader_cmp95_reg == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc163_3_110;
LEGUP_F_main_BB_for_cond92_preheader_preheader_62:
		next_state = LEGUP_F_main_BB_for_cond92_preheader_63;
LEGUP_F_main_BB_for_end214_109:
		next_state = LEGUP_0;
LEGUP_F_main_BB_for_end214_loopexit1_108:
		next_state = LEGUP_F_main_BB_for_end214_109;
LEGUP_F_main_BB_for_end214_loopexit_107:
		next_state = LEGUP_F_main_BB_for_end214_109;
LEGUP_F_main_BB_for_inc163_3_110:
		next_state = LEGUP_F_main_BB_for_inc163_3_111;
LEGUP_F_main_BB_for_inc163_3_111:
		next_state = LEGUP_F_main_BB_for_inc163_3_112;
LEGUP_F_main_BB_for_inc163_3_112:
		next_state = LEGUP_F_main_BB_for_inc166_68;
LEGUP_F_main_BB_for_inc163_us_3_113:
		next_state = LEGUP_F_main_BB_for_inc163_us_3_114;
LEGUP_F_main_BB_for_inc163_us_3_114:
		next_state = LEGUP_F_main_BB_for_inc163_us_3_115;
LEGUP_F_main_BB_for_inc163_us_3_115:
		next_state = LEGUP_F_main_BB_for_inc163_us_3_116;
LEGUP_F_main_BB_for_inc163_us_3_116:
		next_state = LEGUP_F_main_BB_for_inc163_us_3_117;
LEGUP_F_main_BB_for_inc163_us_3_117:
		next_state = LEGUP_F_main_BB_for_inc163_us_3_118;
LEGUP_F_main_BB_for_inc163_us_3_118:
		next_state = LEGUP_F_main_BB_for_inc163_us_3_119;
LEGUP_F_main_BB_for_inc163_us_3_119:
		next_state = LEGUP_F_main_BB_for_inc166_68;
LEGUP_F_main_BB_for_inc166_68:
	if ((fsm_stall == 1'd0) && (main_for_inc166_exitcond12 == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond169_preheader_67;
	else if ((fsm_stall == 1'd0) && (main_for_inc166_exitcond12 == 1'd0))
		next_state = LEGUP_F_main_BB_for_cond92_preheader_63;
LEGUP_F_main_BB_for_inc212_106:
	if ((fsm_stall == 1'd0) && (main_for_inc212_cmp170 == 1'd1))
		next_state = LEGUP_F_main_BB_for_body172_69;
	else if ((fsm_stall == 1'd0) && (main_for_inc212_cmp170 == 1'd0))
		next_state = LEGUP_F_main_BB_for_end214_loopexit1_108;
LEGUP_F_main_BB_for_inc212_loopexit_105:
		next_state = LEGUP_F_main_BB_for_inc212_106;
LEGUP_F_main_BB_for_inc28_i_96:
	if ((fsm_stall == 1'd0) && (main_for_inc28_i_exitcond == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc31_i_97;
	else if ((fsm_stall == 1'd0) && (main_for_inc28_i_exitcond == 1'd0))
		next_state = LEGUP_F_main_BB_for_body11_i_87;
LEGUP_F_main_BB_for_inc31_i_97:
	if ((fsm_stall == 1'd0) && (main_for_inc31_i_exitcond9 == 1'd1))
		next_state = LEGUP_F_main_BB_dijkstra_exit_98;
	else if ((fsm_stall == 1'd0) && (main_for_inc31_i_exitcond9 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body6_i_79;
LEGUP_F_main_BB_for_inc67_15_122:
	if ((fsm_stall == 1'd0) && (main_for_inc67_15_exitcond322 == 1'd1))
		next_state = LEGUP_F_main_BB_for_body75_preheader_123;
	else if ((fsm_stall == 1'd0) && (main_for_inc67_15_exitcond322 == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_124;
LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_124:
		next_state = LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_125;
LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_125:
		next_state = LEGUP_F_main_BB_for_cond58_preheader_28;
LEGUP_F_main_BB_for_inc67_15_storemerge_120:
		next_state = LEGUP_F_main_BB_for_inc67_15_storemerge_121;
LEGUP_F_main_BB_for_inc67_15_storemerge_121:
		next_state = LEGUP_F_main_BB_for_inc67_15_122;
LEGUP_F_main_BB_for_inc_15_128:
	if ((fsm_stall == 1'd0) && (main_for_inc_15_exitcond324 == 1'd1))
		next_state = LEGUP_F_main_BB_for_cond58_preheader_preheader_129;
	else if ((fsm_stall == 1'd0) && (main_for_inc_15_exitcond324 == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_130;
LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_130:
		next_state = LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_131;
LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_131:
		next_state = LEGUP_F_main_BB_for_cond43_preheader_11;
LEGUP_F_main_BB_for_inc_15_storemerge_126:
		next_state = LEGUP_F_main_BB_for_inc_15_storemerge_127;
LEGUP_F_main_BB_for_inc_15_storemerge_127:
		next_state = LEGUP_F_main_BB_for_inc_15_128;
LEGUP_F_main_BB_for_inc_i_i_84:
	if ((fsm_stall == 1'd0) && (main_for_inc_i_i_exitcond2 == 1'd1))
		next_state = LEGUP_F_main_BB_minDistance_exit_i_85;
	else if ((fsm_stall == 1'd0) && (main_for_inc_i_i_exitcond2 == 1'd0))
		next_state = LEGUP_F_main_BB_for_body_i_i_80;
LEGUP_F_main_BB_if_end185_101:
		next_state = LEGUP_F_main_BB_if_end185_102;
LEGUP_F_main_BB_if_end185_102:
	if ((fsm_stall == 1'd0) && (main_if_end185_and192297 == 1'd1))
		next_state = LEGUP_F_main_BB_if_then194_103;
	else if ((fsm_stall == 1'd0) && (main_if_end185_and192297 == 1'd0))
		next_state = LEGUP_F_main_BB_for_end214_loopexit_107;
LEGUP_F_main_BB_if_end185_preheader_100:
		next_state = LEGUP_F_main_BB_if_end185_101;
LEGUP_F_main_BB_if_then194_103:
		next_state = LEGUP_F_main_BB_if_then194_104;
LEGUP_F_main_BB_if_then194_104:
	if ((fsm_stall == 1'd0) && (main_if_then194_cmp182 == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc212_loopexit_105;
	else if ((fsm_stall == 1'd0) && (main_if_then194_cmp182 == 1'd0))
		next_state = LEGUP_F_main_BB_if_end185_101;
LEGUP_F_main_BB_if_then_i_94:
		next_state = LEGUP_F_main_BB_if_then_i_95;
LEGUP_F_main_BB_if_then_i_95:
		next_state = LEGUP_F_main_BB_for_inc28_i_96;
LEGUP_F_main_BB_land_lhs_true16_i_92:
		next_state = LEGUP_F_main_BB_land_lhs_true16_i_93;
LEGUP_F_main_BB_land_lhs_true16_i_93:
	if ((fsm_stall == 1'd0) && (main_land_lhs_true16_i_cmp21_i == 1'd1))
		next_state = LEGUP_F_main_BB_if_then_i_94;
	else if ((fsm_stall == 1'd0) && (main_land_lhs_true16_i_cmp21_i == 1'd0))
		next_state = LEGUP_F_main_BB_for_inc28_i_96;
LEGUP_F_main_BB_land_lhs_true_i_89:
		next_state = LEGUP_F_main_BB_land_lhs_true_i_90;
LEGUP_F_main_BB_land_lhs_true_i_90:
		next_state = LEGUP_F_main_BB_land_lhs_true_i_91;
LEGUP_F_main_BB_land_lhs_true_i_91:
	if ((fsm_stall == 1'd0) && (main_land_lhs_true_i_tobool15_i == 1'd1))
		next_state = LEGUP_F_main_BB_for_inc28_i_96;
	else if ((fsm_stall == 1'd0) && (main_land_lhs_true_i_tobool15_i == 1'd0))
		next_state = LEGUP_F_main_BB_land_lhs_true16_i_92;
LEGUP_F_main_BB_land_lhs_true_i_i_82:
		next_state = LEGUP_F_main_BB_land_lhs_true_i_i_83;
LEGUP_F_main_BB_land_lhs_true_i_i_83:
		next_state = LEGUP_F_main_BB_for_inc_i_i_84;
LEGUP_F_main_BB_minDistance_exit_i_85:
		next_state = LEGUP_F_main_BB_minDistance_exit_i_86;
LEGUP_F_main_BB_minDistance_exit_i_86:
		next_state = LEGUP_F_main_BB_for_body11_i_87;
default:
	next_state = cur_state;
endcase

end
assign fsm_stall = 1'd0;
assign main_entry_0 = 1'd0;
assign main_entry_1 = 1'd0;
assign main_entry_2 = (1'd0 + (4 * 32'd1));
assign main_entry_3 = (1'd0 + (4 * 32'd1));
assign main_entry_4 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_4_reg <= main_entry_4;
	end
end
assign main_entry_5 = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_5_reg <= main_entry_5;
	end
end
assign main_entry_6 = (1'd0 + (4 * 32'd3));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_6_reg <= main_entry_6;
	end
end
assign main_entry_7 = (1'd0 + (4 * 32'd3));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_7_reg <= main_entry_7;
	end
end
assign main_entry_8 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_8_reg <= main_entry_8;
	end
end
assign main_entry_9 = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_9_reg <= main_entry_9;
	end
end
assign main_entry_10 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_10_reg <= main_entry_10;
	end
end
assign main_entry_11 = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_11_reg <= main_entry_11;
	end
end
assign main_entry_12 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_12_reg <= main_entry_12;
	end
end
assign main_entry_13 = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_13_reg <= main_entry_13;
	end
end
assign main_entry_14 = (1'd0 + (4 * 32'd7));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_14_reg <= main_entry_14;
	end
end
assign main_entry_15 = (1'd0 + (4 * 32'd7));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_15_reg <= main_entry_15;
	end
end
assign main_entry_16 = (1'd0 + (4 * 32'd8));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_16_reg <= main_entry_16;
	end
end
assign main_entry_17 = (1'd0 + (4 * 32'd8));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_17_reg <= main_entry_17;
	end
end
assign main_entry_18 = (1'd0 + (4 * 32'd9));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_18_reg <= main_entry_18;
	end
end
assign main_entry_19 = (1'd0 + (4 * 32'd9));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_19_reg <= main_entry_19;
	end
end
assign main_entry_20 = (1'd0 + (4 * 32'd10));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_20_reg <= main_entry_20;
	end
end
assign main_entry_21 = (1'd0 + (4 * 32'd10));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_21_reg <= main_entry_21;
	end
end
assign main_entry_22 = (1'd0 + (4 * 32'd11));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_22_reg <= main_entry_22;
	end
end
assign main_entry_23 = (1'd0 + (4 * 32'd11));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_23_reg <= main_entry_23;
	end
end
assign main_entry_24 = (1'd0 + (4 * 32'd12));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_24_reg <= main_entry_24;
	end
end
assign main_entry_25 = (1'd0 + (4 * 32'd12));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_25_reg <= main_entry_25;
	end
end
assign main_entry_26 = (1'd0 + (4 * 32'd13));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_26_reg <= main_entry_26;
	end
end
assign main_entry_27 = (1'd0 + (4 * 32'd13));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_27_reg <= main_entry_27;
	end
end
assign main_entry_28 = (1'd0 + (4 * 32'd14));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_28_reg <= main_entry_28;
	end
end
assign main_entry_29 = (1'd0 + (4 * 32'd14));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_29_reg <= main_entry_29;
	end
end
assign main_entry_30 = (1'd0 + (4 * 32'd15));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_30_reg <= main_entry_30;
	end
end
assign main_entry_31 = (1'd0 + (4 * 32'd15));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_31_reg <= main_entry_31;
	end
end
assign main_entry_32 = (1'd0 + (4 * 32'd16));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_32_reg <= main_entry_32;
	end
end
assign main_entry_33 = (1'd0 + (4 * 32'd16));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_33_reg <= main_entry_33;
	end
end
assign main_entry_34 = (1'd0 + (4 * 32'd17));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_34_reg <= main_entry_34;
	end
end
assign main_entry_35 = (1'd0 + (4 * 32'd17));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_35_reg <= main_entry_35;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_entry_10) & (fsm_stall == 1'd0))) begin
		main_for_cond43_preheader_36 = 32'd15;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_131) & (fsm_stall == 1'd0))) */ begin
		main_for_cond43_preheader_36 = main_for_inc_15_for_cond43_preheader_crit_edge_pre;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_entry_10) & (fsm_stall == 1'd0))) begin
		main_for_cond43_preheader_36_reg <= main_for_cond43_preheader_36;
	end
	if (((cur_state == LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_131) & (fsm_stall == 1'd0))) begin
		main_for_cond43_preheader_36_reg <= main_for_cond43_preheader_36;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_entry_10) & (fsm_stall == 1'd0))) begin
		main_for_cond43_preheader_37 = 32'd0;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_131) & (fsm_stall == 1'd0))) */ begin
		main_for_cond43_preheader_37 = main_for_cond43_preheader_38_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_entry_10) & (fsm_stall == 1'd0))) begin
		main_for_cond43_preheader_37_reg <= main_for_cond43_preheader_37;
	end
	if (((cur_state == LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_131) & (fsm_stall == 1'd0))) begin
		main_for_cond43_preheader_37_reg <= main_for_cond43_preheader_37;
	end
end
always @(*) begin
		main_for_cond43_preheader_arrayidx49 = (1'd0 + (4 * main_for_cond43_preheader_37_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond43_preheader_11)) begin
		main_for_cond43_preheader_arrayidx49_reg <= main_for_cond43_preheader_arrayidx49;
	end
end
always @(*) begin
		main_for_cond43_preheader_scevgep49 = (1'd0 + (4 * main_for_cond43_preheader_37_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond43_preheader_11)) begin
		main_for_cond43_preheader_scevgep49_reg <= main_for_cond43_preheader_scevgep49;
	end
end
always @(*) begin
		main_for_cond43_preheader_38 = (main_for_cond43_preheader_37_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond43_preheader_11)) begin
		main_for_cond43_preheader_38_reg <= main_for_cond43_preheader_38;
	end
end
always @(*) begin
		main_for_cond43_preheader_Pivot30 = ($signed(main_for_cond43_preheader_36_reg) < $signed({26'd0,main_for_cond43_preheader_Pivot30_op1_temp}));
end
always @(*) begin
		main_NodeBlock27_Pivot28 = ($signed(main_for_cond43_preheader_36_reg) < $signed({26'd0,main_NodeBlock27_Pivot28_op1_temp}));
end
always @(*) begin
		main_NodeBlock25_Pivot26 = ($signed(main_for_cond43_preheader_36_reg) < $signed({26'd0,main_NodeBlock25_Pivot26_op1_temp}));
end
always @(*) begin
		main_NodeBlock23_Pivot24 = ($signed(main_for_cond43_preheader_36_reg) < $signed({26'd0,main_NodeBlock23_Pivot24_op1_temp}));
end
always @(*) begin
		main_LeafBlock21_SwitchLeaf22 = (main_for_cond43_preheader_36_reg == 32'd15);
end
always @(*) begin
		main_NodeBlock19_Pivot20 = ($signed(main_for_cond43_preheader_36_reg) < $signed({26'd0,main_NodeBlock19_Pivot20_op1_temp}));
end
always @(*) begin
		main_NodeBlock19_1 = (main_NodeBlock19_Pivot20 ? 32'd11 : 32'd6);
end
always @(*) begin
		main_NodeBlock17_Pivot18 = ($signed(main_for_cond43_preheader_36_reg) < $signed({26'd0,main_NodeBlock17_Pivot18_op1_temp}));
end
always @(*) begin
		main_NodeBlock15_Pivot16 = ($signed(main_for_cond43_preheader_36_reg) < $signed({26'd0,main_NodeBlock15_Pivot16_op1_temp}));
end
always @(*) begin
		main_NodeBlock15_66 = (main_NodeBlock15_Pivot16 ? 32'd15 : 32'd0);
end
always @(*) begin
		main_NodeBlock13_Pivot14 = ($signed(main_for_cond43_preheader_36_reg) < $signed({26'd0,main_NodeBlock13_Pivot14_op1_temp}));
end
always @(*) begin
		main_NodeBlock13_67 = (main_NodeBlock13_Pivot14 ? 32'd10 : 32'd14);
end
always @(*) begin
		main_NodeBlock11_Pivot12 = ($signed(main_for_cond43_preheader_36_reg) < $signed({27'd0,main_NodeBlock11_Pivot12_op1_temp}));
end
always @(*) begin
		main_NodeBlock9_Pivot10 = ($signed(main_for_cond43_preheader_36_reg) < $signed({27'd0,main_NodeBlock9_Pivot10_op1_temp}));
end
always @(*) begin
		main_NodeBlock7_Pivot8 = ($signed(main_for_cond43_preheader_36_reg) < $signed({27'd0,main_NodeBlock7_Pivot8_op1_temp}));
end
always @(*) begin
		main_NodeBlock7_68 = (main_NodeBlock7_Pivot8 ? 32'd2 : 32'd5);
end
always @(*) begin
		main_NodeBlock5_Pivot6 = ($signed(main_for_cond43_preheader_36_reg) < $signed({27'd0,main_NodeBlock5_Pivot6_op1_temp}));
end
always @(*) begin
		main_NodeBlock5_69 = (main_NodeBlock5_Pivot6 ? 32'd1 : 32'd13);
end
always @(*) begin
		main_NodeBlock3_Pivot4 = ($signed(main_for_cond43_preheader_36_reg) < $signed({28'd0,main_NodeBlock3_Pivot4_op1_temp}));
end
always @(*) begin
		main_NodeBlock1_Pivot2 = ($signed(main_for_cond43_preheader_36_reg) < $signed({28'd0,main_NodeBlock1_Pivot2_op1_temp}));
end
always @(*) begin
		main_NodeBlock1_70 = (main_NodeBlock1_Pivot2 ? 32'd4 : 32'd12);
end
always @(*) begin
		main_NodeBlock_Pivot = ($signed(main_for_cond43_preheader_36_reg) < $signed({29'd0,main_NodeBlock_Pivot_op1_temp}));
end
always @(*) begin
		main_LeafBlock_SwitchLeaf = (main_for_cond43_preheader_36_reg == 32'd0);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_125) & (fsm_stall == 1'd0))) begin
		main_for_cond58_preheader_39 = main_for_inc67_15_for_cond58_preheader_crit_edge_p;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond58_preheader_preheader_129) & (fsm_stall == 1'd0))) */ begin
		main_for_cond58_preheader_39 = 32'd14;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_125) & (fsm_stall == 1'd0))) begin
		main_for_cond58_preheader_39_reg <= main_for_cond58_preheader_39;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond58_preheader_preheader_129) & (fsm_stall == 1'd0))) begin
		main_for_cond58_preheader_39_reg <= main_for_cond58_preheader_39;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_125) & (fsm_stall == 1'd0))) begin
		main_for_cond58_preheader_40 = main_for_cond58_preheader_41_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_cond58_preheader_preheader_129) & (fsm_stall == 1'd0))) */ begin
		main_for_cond58_preheader_40 = 32'd0;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_125) & (fsm_stall == 1'd0))) begin
		main_for_cond58_preheader_40_reg <= main_for_cond58_preheader_40;
	end
	if (((cur_state == LEGUP_F_main_BB_for_cond58_preheader_preheader_129) & (fsm_stall == 1'd0))) begin
		main_for_cond58_preheader_40_reg <= main_for_cond58_preheader_40;
	end
end
always @(*) begin
		main_for_cond58_preheader_arrayidx65 = (1'd0 + (4 * main_for_cond58_preheader_40_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond58_preheader_28)) begin
		main_for_cond58_preheader_arrayidx65_reg <= main_for_cond58_preheader_arrayidx65;
	end
end
always @(*) begin
		main_for_cond58_preheader_scevgep47 = (1'd0 + (4 * main_for_cond58_preheader_40_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond58_preheader_28)) begin
		main_for_cond58_preheader_scevgep47_reg <= main_for_cond58_preheader_scevgep47;
	end
end
always @(*) begin
		main_for_cond58_preheader_41 = (main_for_cond58_preheader_40_reg + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond58_preheader_28)) begin
		main_for_cond58_preheader_41_reg <= main_for_cond58_preheader_41;
	end
end
always @(*) begin
		main_for_cond58_preheader_Pivot65 = ($signed(main_for_cond58_preheader_39_reg) < $signed({26'd0,main_for_cond58_preheader_Pivot65_op1_temp}));
end
always @(*) begin
		main_NodeBlock62_Pivot63 = ($signed(main_for_cond58_preheader_39_reg) < $signed({26'd0,main_NodeBlock62_Pivot63_op1_temp}));
end
always @(*) begin
		main_NodeBlock60_Pivot61 = ($signed(main_for_cond58_preheader_39_reg) < $signed({26'd0,main_NodeBlock60_Pivot61_op1_temp}));
end
always @(*) begin
		main_NodeBlock58_Pivot59 = ($signed(main_for_cond58_preheader_39_reg) < $signed({26'd0,main_NodeBlock58_Pivot59_op1_temp}));
end
always @(*) begin
		main_LeafBlock56_SwitchLeaf57 = (main_for_cond58_preheader_39_reg == 32'd15);
end
always @(*) begin
		main_NodeBlock54_Pivot55 = ($signed(main_for_cond58_preheader_39_reg) < $signed({26'd0,main_NodeBlock54_Pivot55_op1_temp}));
end
always @(*) begin
		main_NodeBlock54_71 = (main_NodeBlock54_Pivot55 ? 32'd11 : 32'd6);
end
always @(*) begin
		main_NodeBlock52_Pivot53 = ($signed(main_for_cond58_preheader_39_reg) < $signed({26'd0,main_NodeBlock52_Pivot53_op1_temp}));
end
always @(*) begin
		main_NodeBlock50_Pivot51 = ($signed(main_for_cond58_preheader_39_reg) < $signed({26'd0,main_NodeBlock50_Pivot51_op1_temp}));
end
always @(*) begin
		main_NodeBlock50_72 = (main_NodeBlock50_Pivot51 ? 32'd15 : 32'd0);
end
always @(*) begin
		main_NodeBlock48_Pivot49 = ($signed(main_for_cond58_preheader_39_reg) < $signed({26'd0,main_NodeBlock48_Pivot49_op1_temp}));
end
always @(*) begin
		main_NodeBlock48_73 = (main_NodeBlock48_Pivot49 ? 32'd10 : 32'd14);
end
always @(*) begin
		main_NodeBlock46_Pivot47 = ($signed(main_for_cond58_preheader_39_reg) < $signed({27'd0,main_NodeBlock46_Pivot47_op1_temp}));
end
always @(*) begin
		main_NodeBlock44_Pivot45 = ($signed(main_for_cond58_preheader_39_reg) < $signed({27'd0,main_NodeBlock44_Pivot45_op1_temp}));
end
always @(*) begin
		main_NodeBlock42_Pivot43 = ($signed(main_for_cond58_preheader_39_reg) < $signed({27'd0,main_NodeBlock42_Pivot43_op1_temp}));
end
always @(*) begin
		main_NodeBlock42_74 = (main_NodeBlock42_Pivot43 ? 32'd2 : 32'd5);
end
always @(*) begin
		main_NodeBlock40_Pivot41 = ($signed(main_for_cond58_preheader_39_reg) < $signed({27'd0,main_NodeBlock40_Pivot41_op1_temp}));
end
always @(*) begin
		main_NodeBlock40_75 = (main_NodeBlock40_Pivot41 ? 32'd1 : 32'd13);
end
always @(*) begin
		main_NodeBlock38_Pivot39 = ($signed(main_for_cond58_preheader_39_reg) < $signed({28'd0,main_NodeBlock38_Pivot39_op1_temp}));
end
always @(*) begin
		main_NodeBlock36_Pivot37 = ($signed(main_for_cond58_preheader_39_reg) < $signed({28'd0,main_NodeBlock36_Pivot37_op1_temp}));
end
always @(*) begin
		main_NodeBlock36_76 = (main_NodeBlock36_Pivot37 ? 32'd4 : 32'd12);
end
always @(*) begin
		main_NodeBlock34_Pivot35 = ($signed(main_for_cond58_preheader_39_reg) < $signed({29'd0,main_NodeBlock34_Pivot35_op1_temp}));
end
always @(*) begin
		main_LeafBlock32_SwitchLeaf33 = (main_for_cond58_preheader_39_reg == 32'd0);
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body75_61) & (fsm_stall == 1'd0)) & (main_for_body75_exitcond59_reg == 1'd0))) begin
		main_for_body75_i_0312 = main_for_body75_42_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_for_body75_preheader_123) & (fsm_stall == 1'd0))) */ begin
		main_for_body75_i_0312 = 32'd0;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body75_61) & (fsm_stall == 1'd0)) & (main_for_body75_exitcond59_reg == 1'd0))) begin
		main_for_body75_i_0312_reg <= main_for_body75_i_0312;
	end
	if (((cur_state == LEGUP_F_main_BB_for_body75_preheader_123) & (fsm_stall == 1'd0))) begin
		main_for_body75_i_0312_reg <= main_for_body75_i_0312;
	end
end
always @(*) begin
		main_for_body75_bit_select7 = main_for_body75_i_0312_reg_width_extended[27:0];
end
always @(*) begin
		main_for_body75_arrayidx76 = (1'd0 + (4 * {27'd0,main_for_body75_i_0312_reg}));
end
always @(*) begin
		main_for_body75_arrayidx77 = (1'd0 + (4 * {27'd0,main_for_body75_i_0312_reg}));
end
always @(*) begin
		main_for_body75_bit_concat23 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat23_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep44 = (1'd0 + (4 * main_for_body75_bit_concat23));
end
always @(*) begin
		main_for_body75_bit_concat22 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat22_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep43 = (1'd0 + (4 * main_for_body75_bit_concat22));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep43_reg <= main_for_body75_scevgep43;
	end
end
always @(*) begin
		main_for_body75_bit_concat21 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat21_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep42 = (1'd0 + (4 * main_for_body75_bit_concat21));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep42_reg <= main_for_body75_scevgep42;
	end
end
always @(*) begin
		main_for_body75_bit_concat20 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat20_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep41 = (1'd0 + (4 * main_for_body75_bit_concat20));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep41_reg <= main_for_body75_scevgep41;
	end
end
always @(*) begin
		main_for_body75_bit_concat19 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat19_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep40 = (1'd0 + (4 * main_for_body75_bit_concat19));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep40_reg <= main_for_body75_scevgep40;
	end
end
always @(*) begin
		main_for_body75_bit_concat18 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat18_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep39 = (1'd0 + (4 * main_for_body75_bit_concat18));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep39_reg <= main_for_body75_scevgep39;
	end
end
always @(*) begin
		main_for_body75_bit_concat17 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat17_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep38 = (1'd0 + (4 * main_for_body75_bit_concat17));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep38_reg <= main_for_body75_scevgep38;
	end
end
always @(*) begin
		main_for_body75_bit_concat16 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat16_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep37 = (1'd0 + (4 * main_for_body75_bit_concat16));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep37_reg <= main_for_body75_scevgep37;
	end
end
always @(*) begin
		main_for_body75_bit_concat15 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat15_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep36 = (1'd0 + (4 * main_for_body75_bit_concat15));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep36_reg <= main_for_body75_scevgep36;
	end
end
always @(*) begin
		main_for_body75_bit_concat14 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat14_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep35 = (1'd0 + (4 * main_for_body75_bit_concat14));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep35_reg <= main_for_body75_scevgep35;
	end
end
always @(*) begin
		main_for_body75_bit_concat13 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat13_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep34 = (1'd0 + (4 * main_for_body75_bit_concat13));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep34_reg <= main_for_body75_scevgep34;
	end
end
always @(*) begin
		main_for_body75_bit_concat12 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat12_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep33 = (1'd0 + (4 * main_for_body75_bit_concat12));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep33_reg <= main_for_body75_scevgep33;
	end
end
always @(*) begin
		main_for_body75_bit_concat11 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat11_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep32 = (1'd0 + (4 * main_for_body75_bit_concat11));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep32_reg <= main_for_body75_scevgep32;
	end
end
always @(*) begin
		main_for_body75_bit_concat10 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat10_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep31 = (1'd0 + (4 * main_for_body75_bit_concat10));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep31_reg <= main_for_body75_scevgep31;
	end
end
always @(*) begin
		main_for_body75_bit_concat9 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat9_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep30 = (1'd0 + (4 * main_for_body75_bit_concat9));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep30_reg <= main_for_body75_scevgep30;
	end
end
always @(*) begin
		main_for_body75_bit_concat8 = {main_for_body75_bit_select7[27:0], main_for_body75_bit_concat8_bit_select_operand_2[3:0]};
end
always @(*) begin
		main_for_body75_scevgep29 = (1'd0 + (4 * main_for_body75_bit_concat8));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_scevgep29_reg <= main_for_body75_scevgep29;
	end
end
always @(*) begin
		main_for_body75_42 = ({1'd0,main_for_body75_i_0312_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_42_reg <= main_for_body75_42;
	end
end
always @(*) begin
		main_for_body75_exitcond59 = (main_for_body75_42 == 32'd16);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_for_body75_exitcond59_reg <= main_for_body75_exitcond59;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond92_preheader_preheader_62) & (fsm_stall == 1'd0))) begin
		main_for_cond92_preheader_43 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc166_68) & (fsm_stall == 1'd0)) & (main_for_inc166_exitcond12 == 1'd0))) */ begin
		main_for_cond92_preheader_43 = main_for_inc166_49;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond92_preheader_preheader_62) & (fsm_stall == 1'd0))) begin
		main_for_cond92_preheader_43_reg <= main_for_cond92_preheader_43;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc166_68) & (fsm_stall == 1'd0)) & (main_for_inc166_exitcond12 == 1'd0))) begin
		main_for_cond92_preheader_43_reg <= main_for_cond92_preheader_43;
	end
end
always @(*) begin
		main_for_cond92_preheader_bit_select5 = main_for_cond92_preheader_43_reg_width_extended[29:0];
end
always @(*) begin
		main_for_cond92_preheader_bit_select3 = main_for_cond92_preheader_43_reg_width_extended[25:0];
end
always @(*) begin
		main_for_cond92_preheader_bit_concat6 = {main_for_cond92_preheader_bit_select5[29:0], main_for_cond92_preheader_bit_concat6_bit_select_operand_2[1:0]};
end
always @(*) begin
		main_for_cond92_preheader_bit_concat4 = {main_for_cond92_preheader_bit_select3[25:0], main_for_cond92_preheader_bit_concat4_bit_select_operand_2[5:0]};
end
always @(*) begin
		main_for_cond92_preheader_sr_add = (main_for_cond92_preheader_bit_concat6 + main_for_cond92_preheader_bit_concat4);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_63)) begin
		main_for_cond92_preheader_sr_add_reg <= main_for_cond92_preheader_sr_add;
	end
end
always @(*) begin
		main_for_cond92_preheader_bit_select1 = main_for_cond92_preheader_sr_add[31:1];
end
always @(*) begin
		main_for_cond92_preheader_44 = (main_for_cond92_preheader_sr_add + 32'd16);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_63)) begin
		main_for_cond92_preheader_44_reg <= main_for_cond92_preheader_44;
	end
end
always @(*) begin
		main_for_cond92_preheader_scevgep27 = (1'd0 + (4 * main_for_cond92_preheader_44_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_64)) begin
		main_for_cond92_preheader_scevgep27_reg <= main_for_cond92_preheader_scevgep27;
	end
end
always @(*) begin
		main_for_cond92_preheader_bit_concat2 = {main_for_cond92_preheader_bit_select1[30:0], main_for_cond92_preheader_bit_concat2_bit_select_operand_2};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_63)) begin
		main_for_cond92_preheader_bit_concat2_reg <= main_for_cond92_preheader_bit_concat2;
	end
end
always @(*) begin
		main_for_cond92_preheader_scevgep26 = (1'd0 + (4 * main_for_cond92_preheader_bit_concat2_reg));
end
always @(*) begin
		main_for_cond92_preheader_45 = (main_for_cond92_preheader_sr_add + 32'd33);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_63)) begin
		main_for_cond92_preheader_45_reg <= main_for_cond92_preheader_45;
	end
end
always @(*) begin
		main_for_cond92_preheader_scevgep25 = (1'd0 + (4 * main_for_cond92_preheader_45_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_64)) begin
		main_for_cond92_preheader_scevgep25_reg <= main_for_cond92_preheader_scevgep25;
	end
end
always @(*) begin
		main_for_cond92_preheader_46 = (main_for_cond92_preheader_sr_add + 32'd50);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_63)) begin
		main_for_cond92_preheader_46_reg <= main_for_cond92_preheader_46;
	end
end
always @(*) begin
		main_for_cond92_preheader_scevgep23 = (1'd0 + (4 * main_for_cond92_preheader_46_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_64)) begin
		main_for_cond92_preheader_scevgep23_reg <= main_for_cond92_preheader_scevgep23;
	end
end
always @(*) begin
		main_for_cond92_preheader_47 = (main_for_cond92_preheader_sr_add + 32'd18);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_63)) begin
		main_for_cond92_preheader_47_reg <= main_for_cond92_preheader_47;
	end
end
always @(*) begin
		main_for_cond92_preheader_scevgep22 = (1'd0 + (4 * main_for_cond92_preheader_47_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_64)) begin
		main_for_cond92_preheader_scevgep22_reg <= main_for_cond92_preheader_scevgep22;
	end
end
always @(*) begin
		main_for_cond92_preheader_48 = (main_for_cond92_preheader_sr_add + 32'd35);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_63)) begin
		main_for_cond92_preheader_48_reg <= main_for_cond92_preheader_48;
	end
end
always @(*) begin
		main_for_cond92_preheader_scevgep20 = (1'd0 + (4 * main_for_cond92_preheader_48_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_64)) begin
		main_for_cond92_preheader_scevgep20_reg <= main_for_cond92_preheader_scevgep20;
	end
end
always @(*) begin
		main_for_cond92_preheader_cmp95 = ($signed({28'd0,main_for_cond92_preheader_cmp95_op0_temp}) < $signed({28'd0,main_for_cond92_preheader_cmp95_op1_temp}));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_63)) begin
		main_for_cond92_preheader_cmp95_reg <= main_for_cond92_preheader_cmp95;
	end
end
assign main_for_cond169_preheader_arrayidx1_i = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_i_reg <= main_for_cond169_preheader_arrayidx1_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_i = 1'd0;
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_i_reg <= main_for_cond169_preheader_arrayidx2_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_1_i = (1'd0 + (4 * 32'd1));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_1_i_reg <= main_for_cond169_preheader_arrayidx1_1_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_1_i = (1'd0 + (4 * 32'd1));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_1_i_reg <= main_for_cond169_preheader_arrayidx2_1_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_2_i = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_2_i_reg <= main_for_cond169_preheader_arrayidx1_2_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_2_i = (1'd0 + (4 * 32'd2));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_2_i_reg <= main_for_cond169_preheader_arrayidx2_2_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_3_i = (1'd0 + (4 * 32'd3));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_3_i_reg <= main_for_cond169_preheader_arrayidx1_3_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_3_i = (1'd0 + (4 * 32'd3));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_3_i_reg <= main_for_cond169_preheader_arrayidx2_3_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_4_i = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_4_i_reg <= main_for_cond169_preheader_arrayidx1_4_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_4_i = (1'd0 + (4 * 32'd4));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_4_i_reg <= main_for_cond169_preheader_arrayidx2_4_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_5_i = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_5_i_reg <= main_for_cond169_preheader_arrayidx1_5_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_5_i = (1'd0 + (4 * 32'd5));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_5_i_reg <= main_for_cond169_preheader_arrayidx2_5_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_6_i = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_6_i_reg <= main_for_cond169_preheader_arrayidx1_6_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_6_i = (1'd0 + (4 * 32'd6));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_6_i_reg <= main_for_cond169_preheader_arrayidx2_6_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_7_i = (1'd0 + (4 * 32'd7));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_7_i_reg <= main_for_cond169_preheader_arrayidx1_7_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_7_i = (1'd0 + (4 * 32'd7));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_7_i_reg <= main_for_cond169_preheader_arrayidx2_7_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_8_i = (1'd0 + (4 * 32'd8));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_8_i_reg <= main_for_cond169_preheader_arrayidx1_8_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_8_i = (1'd0 + (4 * 32'd8));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_8_i_reg <= main_for_cond169_preheader_arrayidx2_8_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_9_i = (1'd0 + (4 * 32'd9));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_9_i_reg <= main_for_cond169_preheader_arrayidx1_9_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_9_i = (1'd0 + (4 * 32'd9));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_9_i_reg <= main_for_cond169_preheader_arrayidx2_9_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_10_i = (1'd0 + (4 * 32'd10));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_10_i_reg <= main_for_cond169_preheader_arrayidx1_10_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_10_i = (1'd0 + (4 * 32'd10));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_10_i_reg <= main_for_cond169_preheader_arrayidx2_10_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_11_i = (1'd0 + (4 * 32'd11));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_11_i_reg <= main_for_cond169_preheader_arrayidx1_11_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_11_i = (1'd0 + (4 * 32'd11));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_11_i_reg <= main_for_cond169_preheader_arrayidx2_11_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_12_i = (1'd0 + (4 * 32'd12));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_12_i_reg <= main_for_cond169_preheader_arrayidx1_12_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_12_i = (1'd0 + (4 * 32'd12));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_12_i_reg <= main_for_cond169_preheader_arrayidx2_12_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_13_i = (1'd0 + (4 * 32'd13));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_13_i_reg <= main_for_cond169_preheader_arrayidx1_13_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_13_i = (1'd0 + (4 * 32'd13));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_13_i_reg <= main_for_cond169_preheader_arrayidx2_13_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_14_i = (1'd0 + (4 * 32'd14));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_14_i_reg <= main_for_cond169_preheader_arrayidx1_14_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_14_i = (1'd0 + (4 * 32'd14));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_14_i_reg <= main_for_cond169_preheader_arrayidx2_14_i;
	end
end
assign main_for_cond169_preheader_arrayidx1_15_i = (1'd0 + (4 * 32'd15));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx1_15_i_reg <= main_for_cond169_preheader_arrayidx1_15_i;
	end
end
assign main_for_cond169_preheader_arrayidx2_15_i = (1'd0 + (4 * 32'd15));
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67)) begin
		main_for_cond169_preheader_arrayidx2_15_i_reg <= main_for_cond169_preheader_arrayidx2_15_i;
	end
end
always @(*) begin
		main_for_inc166_49 = ({1'd0,main_for_cond92_preheader_43_reg} + 32'd1);
end
always @(*) begin
		main_for_inc166_exitcond12 = (main_for_inc166_49 == 32'd4);
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67) & (fsm_stall == 1'd0))) begin
		main_for_body172_i_2307 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc212_106) & (fsm_stall == 1'd0)) & (main_for_inc212_cmp170 == 1'd1))) */ begin
		main_for_body172_i_2307 = main_for_body172_inc213_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_cond169_preheader_67) & (fsm_stall == 1'd0))) begin
		main_for_body172_i_2307_reg <= main_for_body172_i_2307;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc212_106) & (fsm_stall == 1'd0)) & (main_for_inc212_cmp170 == 1'd1))) begin
		main_for_body172_i_2307_reg <= main_for_body172_i_2307;
	end
end
always @(*) begin
		main_for_body172_arrayidx173 = (1'd0 + (4 * {27'd0,main_for_body172_i_2307_reg}));
end
always @(*) begin
		main_for_body172_arrayidx174 = (1'd0 + (4 * {27'd0,main_for_body172_i_2307_reg}));
end
always @(*) begin
		main_for_body172_inc213 = ({1'd0,main_for_body172_i_2307_reg} + 32'd1);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_for_body172_inc213_reg <= main_for_body172_inc213;
	end
end
always @(*) begin
		main_for_body172_50 = main_entry_vla39295_out_a;
end
always @(*) begin
		main_for_body172_51 = main_entry_vla40296_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_for_body172_51_reg <= main_for_body172_51;
	end
end
always @(*) begin
		main_for_body172_arrayidx_i = (1'd0 + (4 * main_for_body172_50));
end
always @(*) begin
		main_for_body172_arrayidx3_i = (1'd0 + (4 * main_for_body172_50));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_for_body172_arrayidx3_i_reg <= main_for_body172_arrayidx3_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body172_78) & (fsm_stall == 1'd0))) begin
		main_for_body6_i_count_056_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc31_i_97) & (fsm_stall == 1'd0)) & (main_for_inc31_i_exitcond9 == 1'd0))) */ begin
		main_for_body6_i_count_056_i = main_for_inc31_i_62;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body172_78) & (fsm_stall == 1'd0))) begin
		main_for_body6_i_count_056_i_reg <= main_for_body6_i_count_056_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc31_i_97) & (fsm_stall == 1'd0)) & (main_for_inc31_i_exitcond9 == 1'd0))) begin
		main_for_body6_i_count_056_i_reg <= main_for_body6_i_count_056_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_79) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_52 = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_84) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond2 == 1'd0))) */ begin
		main_for_body_i_i_52 = main_for_inc_i_i_55;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_79) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_52_reg <= main_for_body_i_i_52;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_84) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond2 == 1'd0))) begin
		main_for_body_i_i_52_reg <= main_for_body_i_i_52;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_79) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_index_012_i_i = 0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_84) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond2 == 1'd0))) */ begin
		main_for_body_i_i_min_index_012_i_i = main_for_inc_i_i_min_index_1_i_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_79) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_index_012_i_i_reg <= main_for_body_i_i_min_index_012_i_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_84) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond2 == 1'd0))) begin
		main_for_body_i_i_min_index_012_i_i_reg <= main_for_body_i_i_min_index_012_i_i;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_79) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_011_i_i = 32'd2147483647;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_84) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond2 == 1'd0))) */ begin
		main_for_body_i_i_min_011_i_i = main_for_inc_i_i_min_1_i_i_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_for_body6_i_79) & (fsm_stall == 1'd0))) begin
		main_for_body_i_i_min_011_i_i_reg <= main_for_body_i_i_min_011_i_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc_i_i_84) & (fsm_stall == 1'd0)) & (main_for_inc_i_i_exitcond2 == 1'd0))) begin
		main_for_body_i_i_min_011_i_i_reg <= main_for_body_i_i_min_011_i_i;
	end
end
always @(*) begin
		main_for_body_i_i_arrayidx_i_i = (1'd0 + (4 * main_for_body_i_i_52_reg));
end
always @(*) begin
		main_for_body_i_i_53 = main_entry_sptSet_i_out_a;
end
always @(*) begin
		main_for_body_i_i_cmp1_i_i = (main_for_body_i_i_53 == 32'd0);
end
always @(*) begin
		main_land_lhs_true_i_i_arrayidx2_i_i = (1'd0 + (4 * main_for_body_i_i_52_reg));
end
always @(*) begin
		main_land_lhs_true_i_i_54 = main_entry_dist_i_out_b;
end
always @(*) begin
		main_land_lhs_true_i_i_cmp3_i_i = ($signed(main_land_lhs_true_i_i_54) > $signed(main_for_body_i_i_min_011_i_i_reg));
end
always @(*) begin
		main_land_lhs_true_i_i_min_0_i_i = (main_land_lhs_true_i_i_cmp3_i_i ? main_for_body_i_i_min_011_i_i_reg : main_land_lhs_true_i_i_54);
end
always @(*) begin
		main_land_lhs_true_i_i_min_index_0_v_0_i_i = (main_land_lhs_true_i_i_cmp3_i_i ? main_for_body_i_i_min_index_012_i_i_reg : main_for_body_i_i_52_reg);
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_81) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_1_i_i = main_for_body_i_i_min_011_i_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_83) & (fsm_stall == 1'd0))) */ begin
		main_for_inc_i_i_min_1_i_i = main_land_lhs_true_i_i_min_0_i_i;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_81) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_1_i_i_reg <= main_for_inc_i_i_min_1_i_i;
	end
	if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_83) & (fsm_stall == 1'd0))) begin
		main_for_inc_i_i_min_1_i_i_reg <= main_for_inc_i_i_min_1_i_i;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_81) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_index_1_i_i = main_for_body_i_i_min_index_012_i_i_reg;
	end
	else /* if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_83) & (fsm_stall == 1'd0))) */ begin
		main_for_inc_i_i_min_index_1_i_i = main_land_lhs_true_i_i_min_index_0_v_0_i_i;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_for_body_i_i_81) & (fsm_stall == 1'd0)) & (main_for_body_i_i_cmp1_i_i == 1'd0))) begin
		main_for_inc_i_i_min_index_1_i_i_reg <= main_for_inc_i_i_min_index_1_i_i;
	end
	if (((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_83) & (fsm_stall == 1'd0))) begin
		main_for_inc_i_i_min_index_1_i_i_reg <= main_for_inc_i_i_min_index_1_i_i;
	end
end
always @(*) begin
		main_for_inc_i_i_bit_select = main_for_inc_i_i_min_index_1_i_i_reg[27:0];
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc_i_i_84)) begin
		main_for_inc_i_i_bit_select_reg <= main_for_inc_i_i_bit_select;
	end
end
always @(*) begin
		main_for_inc_i_i_55 = (main_for_body_i_i_52_reg + 32'd1);
end
always @(*) begin
		main_for_inc_i_i_exitcond2 = (main_for_inc_i_i_55 == 32'd16);
end
always @(*) begin
		main_minDistance_exit_i_arrayidx8_i = (1'd0 + (4 * main_for_inc_i_i_min_index_1_i_i_reg));
end
always @(*) begin
		main_minDistance_exit_i_arrayidx17_i = (1'd0 + (4 * main_for_inc_i_i_min_index_1_i_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_85)) begin
		main_minDistance_exit_i_arrayidx17_i_reg <= main_minDistance_exit_i_arrayidx17_i;
	end
end
always @(*) begin
		main_minDistance_exit_i_bit_concat = {main_for_inc_i_i_bit_select_reg[27:0], main_minDistance_exit_i_bit_concat_bit_select_operand_2[3:0]};
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_85)) begin
		main_minDistance_exit_i_bit_concat_reg <= main_minDistance_exit_i_bit_concat;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_minDistance_exit_i_86) & (fsm_stall == 1'd0))) begin
		main_for_body11_i_v_055_i = 32'd0;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_for_inc28_i_96) & (fsm_stall == 1'd0)) & (main_for_inc28_i_exitcond == 1'd0))) */ begin
		main_for_body11_i_v_055_i = main_for_inc28_i_61;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_minDistance_exit_i_86) & (fsm_stall == 1'd0))) begin
		main_for_body11_i_v_055_i_reg <= main_for_body11_i_v_055_i;
	end
	if ((((cur_state == LEGUP_F_main_BB_for_inc28_i_96) & (fsm_stall == 1'd0)) & (main_for_inc28_i_exitcond == 1'd0))) begin
		main_for_body11_i_v_055_i_reg <= main_for_body11_i_v_055_i;
	end
end
always @(*) begin
		main_for_body11_i_arrayidx12_i = (1'd0 + (4 * main_for_body11_i_v_055_i_reg));
end
always @(*) begin
		main_for_body11_i_arrayidx20_i = (1'd0 + (4 * main_for_body11_i_v_055_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body11_i_87)) begin
		main_for_body11_i_arrayidx20_i_reg <= main_for_body11_i_arrayidx20_i;
	end
end
always @(*) begin
		main_for_body11_i_arrayidx22_i = (1'd0 + (4 * main_for_body11_i_v_055_i_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_body11_i_87)) begin
		main_for_body11_i_arrayidx22_i_reg <= main_for_body11_i_arrayidx22_i;
	end
end
always @(*) begin
		main_for_body11_i_56 = main_entry_sptSet_i_out_a;
end
always @(*) begin
		main_for_body11_i_tobool_i = (main_for_body11_i_56 == 32'd0);
end
always @(*) begin
		main_land_lhs_true_i_57 = (main_minDistance_exit_i_bit_concat_reg + main_for_body11_i_v_055_i_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_89)) begin
		main_land_lhs_true_i_57_reg <= main_land_lhs_true_i_57;
	end
end
always @(*) begin
		main_land_lhs_true_i_scevgep = (1'd0 + (4 * main_land_lhs_true_i_57_reg));
end
always @(*) begin
		main_land_lhs_true_i_58 = main_entry_m1_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_91)) begin
		main_land_lhs_true_i_58_reg <= main_land_lhs_true_i_58;
	end
end
always @(*) begin
		main_land_lhs_true_i_tobool15_i = (main_land_lhs_true_i_58 == 32'd0);
end
always @(*) begin
		main_land_lhs_true16_i_59 = main_entry_dist_i_out_a;
end
always @(*) begin
		main_land_lhs_true16_i_add_i = (main_land_lhs_true16_i_59 + main_land_lhs_true_i_58_reg);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true16_i_93)) begin
		main_land_lhs_true16_i_add_i_reg <= main_land_lhs_true16_i_add_i;
	end
end
always @(*) begin
		main_land_lhs_true16_i_60 = main_entry_dist_i_out_b;
end
always @(*) begin
		main_land_lhs_true16_i_cmp21_i = ($signed(main_land_lhs_true16_i_add_i) < $signed(main_land_lhs_true16_i_60));
end
always @(*) begin
		main_for_inc28_i_61 = (main_for_body11_i_v_055_i_reg + 32'd1);
end
always @(*) begin
		main_for_inc28_i_exitcond = (main_for_inc28_i_61 == 32'd16);
end
always @(*) begin
		main_for_inc31_i_62 = (main_for_body6_i_count_056_i_reg + 32'd1);
end
always @(*) begin
		main_for_inc31_i_exitcond9 = (main_for_inc31_i_62 == 32'd15);
end
always @(*) begin
		main_dijkstra_exit_arrayidx181303 = (1'd0 + (4 * main_for_body172_51_reg));
end
always @(*) begin
		main_dijkstra_exit_63 = main_entry_parent_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_dijkstra_exit_99)) begin
		main_dijkstra_exit_63_reg <= main_dijkstra_exit_63;
	end
end
always @(*) begin
		main_dijkstra_exit_cmp182304 = (main_dijkstra_exit_63 == $signed(-32'd1));
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_end185_preheader_100) & (fsm_stall == 1'd0))) begin
		main_if_end185_64 = main_dijkstra_exit_63_reg;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_if_then194_104) & (fsm_stall == 1'd0)) & (main_if_then194_cmp182 == 1'd0))) */ begin
		main_if_end185_64 = main_if_then194_67;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_end185_preheader_100) & (fsm_stall == 1'd0))) begin
		main_if_end185_64_reg <= main_if_end185_64;
	end
	if ((((cur_state == LEGUP_F_main_BB_if_then194_104) & (fsm_stall == 1'd0)) & (main_if_then194_cmp182 == 1'd0))) begin
		main_if_end185_64_reg <= main_if_end185_64;
	end
end
always @(*) begin
	if (((cur_state == LEGUP_F_main_BB_if_end185_preheader_100) & (fsm_stall == 1'd0))) begin
		main_if_end185_origem_1306 = main_for_body172_51_reg;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_if_then194_104) & (fsm_stall == 1'd0)) & (main_if_then194_cmp182 == 1'd0))) */ begin
		main_if_end185_origem_1306 = main_if_end185_64_reg;
	end
end
always @(posedge clk) begin
	if (((cur_state == LEGUP_F_main_BB_if_end185_preheader_100) & (fsm_stall == 1'd0))) begin
		main_if_end185_origem_1306_reg <= main_if_end185_origem_1306;
	end
	if ((((cur_state == LEGUP_F_main_BB_if_then194_104) & (fsm_stall == 1'd0)) & (main_if_then194_cmp182 == 1'd0))) begin
		main_if_end185_origem_1306_reg <= main_if_end185_origem_1306;
	end
end
always @(*) begin
		main_if_end185_arrayidx186 = (1'd0 + (4 * main_if_end185_64_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end185_101)) begin
		main_if_end185_arrayidx186_reg <= main_if_end185_arrayidx186;
	end
end
always @(*) begin
		main_if_end185_65 = main_entry_indice_s_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end185_102)) begin
		main_if_end185_65_reg <= main_if_end185_65;
	end
end
always @(*) begin
		main_if_end185_cmp187 = ($signed(main_if_end185_65) < $signed({27'd0,main_if_end185_cmp187_op1_temp}));
end
always @(*) begin
		main_if_end185_arrayidx189 = (1'd0 + (4 * main_if_end185_origem_1306_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end185_101)) begin
		main_if_end185_arrayidx189_reg <= main_if_end185_arrayidx189;
	end
end
always @(*) begin
		main_if_end185_66 = main_entry_indice_e_out_a;
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_if_end185_102)) begin
		main_if_end185_66_reg <= main_if_end185_66;
	end
end
always @(*) begin
		main_if_end185_cmp190 = ($signed(main_if_end185_66) < $signed({27'd0,main_if_end185_cmp190_op1_temp}));
end
always @(*) begin
		main_if_end185_and192297 = (main_if_end185_cmp187 & main_if_end185_cmp190);
end
always @(*) begin
		main_if_then194_add202 = (main_if_end185_66_reg + 32'd1);
end
always @(*) begin
		main_if_then194_add204 = (main_if_end185_65_reg + 32'd1);
end
always @(*) begin
		main_if_then194_arrayidx181 = (1'd0 + (4 * main_if_end185_64_reg));
end
always @(*) begin
		main_if_then194_67 = main_entry_parent_out_a;
end
always @(*) begin
		main_if_then194_cmp182 = (main_if_then194_67 == $signed(-32'd1));
end
always @(*) begin
		main_for_inc212_cmp170 = ($signed({25'd0,main_for_inc212_cmp170_op0_temp}) < $signed({25'd0,main_for_inc212_cmp170_op1_temp}));
end
always @(*) begin
		main_for_inc163_us_3_68 = (main_for_cond92_preheader_sr_add_reg + 32'd81);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_for_inc163_us_3_68_reg <= main_for_inc163_us_3_68;
	end
end
always @(*) begin
		main_for_inc163_us_3_scevgep24 = (1'd0 + (4 * main_for_inc163_us_3_68_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_for_inc163_us_3_scevgep24_reg <= main_for_inc163_us_3_scevgep24;
	end
end
always @(*) begin
		main_for_inc163_us_3_69 = (main_for_cond92_preheader_sr_add_reg + 32'd98);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_for_inc163_us_3_69_reg <= main_for_inc163_us_3_69;
	end
end
always @(*) begin
		main_for_inc163_us_3_scevgep21 = (1'd0 + (4 * main_for_inc163_us_3_69_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_for_inc163_us_3_scevgep21_reg <= main_for_inc163_us_3_scevgep21;
	end
end
always @(*) begin
		main_for_inc163_us_3_70 = (main_for_cond92_preheader_sr_add_reg + 32'd115);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_for_inc163_us_3_70_reg <= main_for_inc163_us_3_70;
	end
end
always @(*) begin
		main_for_inc163_us_3_scevgep19 = (1'd0 + (4 * main_for_inc163_us_3_70_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_for_inc163_us_3_scevgep19_reg <= main_for_inc163_us_3_scevgep19;
	end
end
always @(*) begin
		main_for_inc163_us_3_71 = (main_for_cond92_preheader_sr_add_reg + 32'd55);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_for_inc163_us_3_71_reg <= main_for_inc163_us_3_71;
	end
end
always @(*) begin
		main_for_inc163_us_3_scevgep18 = (1'd0 + (4 * main_for_inc163_us_3_71_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_for_inc163_us_3_scevgep18_reg <= main_for_inc163_us_3_scevgep18;
	end
end
always @(*) begin
		main_for_inc163_us_3_72 = (main_for_cond92_preheader_sr_add_reg + 32'd38);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_for_inc163_us_3_72_reg <= main_for_inc163_us_3_72;
	end
end
always @(*) begin
		main_for_inc163_us_3_scevgep17 = (1'd0 + (4 * main_for_inc163_us_3_72_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_for_inc163_us_3_scevgep17_reg <= main_for_inc163_us_3_scevgep17;
	end
end
always @(*) begin
		main_for_inc163_us_3_73 = (main_for_cond92_preheader_sr_add_reg + 32'd21);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_for_inc163_us_3_73_reg <= main_for_inc163_us_3_73;
	end
end
always @(*) begin
		main_for_inc163_us_3_scevgep16 = (1'd0 + (4 * main_for_inc163_us_3_73_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_for_inc163_us_3_scevgep16_reg <= main_for_inc163_us_3_scevgep16;
	end
end
always @(*) begin
		main_for_inc163_us_3_74 = (main_for_cond92_preheader_sr_add_reg + 32'd64);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_for_inc163_us_3_74_reg <= main_for_inc163_us_3_74;
	end
end
always @(*) begin
		main_for_inc163_us_3_scevgep15 = (1'd0 + (4 * main_for_inc163_us_3_74_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_for_inc163_us_3_scevgep15_reg <= main_for_inc163_us_3_scevgep15;
	end
end
always @(*) begin
		main_for_inc163_us_3_75 = (main_for_cond92_preheader_sr_add_reg + 32'd4);
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_for_inc163_us_3_75_reg <= main_for_inc163_us_3_75;
	end
end
always @(*) begin
		main_for_inc163_us_3_scevgep14 = (1'd0 + (4 * main_for_inc163_us_3_75_reg));
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_for_inc163_us_3_scevgep14_reg <= main_for_inc163_us_3_scevgep14;
	end
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock58_31) & (fsm_stall == 1'd0)) & (main_NodeBlock58_Pivot59 == 1'd1))) begin
		main_for_inc67_15_storemerge_storemerge52 = 32'd7;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock56_32) & (fsm_stall == 1'd0)) & (main_LeafBlock56_SwitchLeaf57 == 1'd1))) begin
		main_for_inc67_15_storemerge_storemerge52 = 32'd3;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock54_33) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52 = main_NodeBlock54_71;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock50_35) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52 = main_NodeBlock50_72;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock48_36) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52 = main_NodeBlock48_73;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock42_39) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52 = {1'd0,main_NodeBlock42_74};
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock40_40) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52 = main_NodeBlock40_75;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock36_42) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52 = main_NodeBlock36_76;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock34_43) & (fsm_stall == 1'd0)) & (main_NodeBlock34_Pivot35 == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52 = 32'd9;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_LeafBlock32_44) & (fsm_stall == 1'd0)) & (main_LeafBlock32_SwitchLeaf33 == 1'd1))) */ begin
		main_for_inc67_15_storemerge_storemerge52 = 32'd8;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock58_31) & (fsm_stall == 1'd0)) & (main_NodeBlock58_Pivot59 == 1'd1))) begin
		main_for_inc67_15_storemerge_storemerge52_reg <= main_for_inc67_15_storemerge_storemerge52;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock56_32) & (fsm_stall == 1'd0)) & (main_LeafBlock56_SwitchLeaf57 == 1'd1))) begin
		main_for_inc67_15_storemerge_storemerge52_reg <= main_for_inc67_15_storemerge_storemerge52;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock54_33) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52_reg <= main_for_inc67_15_storemerge_storemerge52;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock50_35) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52_reg <= main_for_inc67_15_storemerge_storemerge52;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock48_36) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52_reg <= main_for_inc67_15_storemerge_storemerge52;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock42_39) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52_reg <= main_for_inc67_15_storemerge_storemerge52;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock40_40) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52_reg <= main_for_inc67_15_storemerge_storemerge52;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock36_42) & (fsm_stall == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52_reg <= main_for_inc67_15_storemerge_storemerge52;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock34_43) & (fsm_stall == 1'd0)) & (main_NodeBlock34_Pivot35 == 1'd0))) begin
		main_for_inc67_15_storemerge_storemerge52_reg <= main_for_inc67_15_storemerge_storemerge52;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock32_44) & (fsm_stall == 1'd0)) & (main_LeafBlock32_SwitchLeaf33 == 1'd1))) begin
		main_for_inc67_15_storemerge_storemerge52_reg <= main_for_inc67_15_storemerge_storemerge52;
	end
end
always @(*) begin
		main_for_inc67_15_exitcond322 = (main_for_cond58_preheader_40_reg == 32'd18);
end
always @(*) begin
		main_for_inc67_15_for_cond58_preheader_crit_edge_p = main_entry_vla12943_out_a;
end
always @(*) begin
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock23_14) & (fsm_stall == 1'd0)) & (main_NodeBlock23_Pivot24 == 1'd1))) begin
		main_for_inc_15_storemerge_storemerge = 32'd7;
	end
	else if ((((cur_state == LEGUP_F_main_BB_LeafBlock21_15) & (fsm_stall == 1'd0)) & (main_LeafBlock21_SwitchLeaf22 == 1'd1))) begin
		main_for_inc_15_storemerge_storemerge = 32'd3;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock19_16) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge = main_NodeBlock19_1;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock15_18) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge = main_NodeBlock15_66;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock13_19) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge = main_NodeBlock13_67;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock7_22) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge = {1'd0,main_NodeBlock7_68};
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock5_23) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge = main_NodeBlock5_69;
	end
	else if (((cur_state == LEGUP_F_main_BB_NodeBlock1_25) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge = main_NodeBlock1_70;
	end
	else if ((((cur_state == LEGUP_F_main_BB_NodeBlock_26) & (fsm_stall == 1'd0)) & (main_NodeBlock_Pivot == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge = 32'd9;
	end
	else /* if ((((cur_state == LEGUP_F_main_BB_LeafBlock_27) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) */ begin
		main_for_inc_15_storemerge_storemerge = 32'd8;
	end
end
always @(posedge clk) begin
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock23_14) & (fsm_stall == 1'd0)) & (main_NodeBlock23_Pivot24 == 1'd1))) begin
		main_for_inc_15_storemerge_storemerge_reg <= main_for_inc_15_storemerge_storemerge;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock21_15) & (fsm_stall == 1'd0)) & (main_LeafBlock21_SwitchLeaf22 == 1'd1))) begin
		main_for_inc_15_storemerge_storemerge_reg <= main_for_inc_15_storemerge_storemerge;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock19_16) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge_reg <= main_for_inc_15_storemerge_storemerge;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock15_18) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge_reg <= main_for_inc_15_storemerge_storemerge;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock13_19) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge_reg <= main_for_inc_15_storemerge_storemerge;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock7_22) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge_reg <= main_for_inc_15_storemerge_storemerge;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock5_23) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge_reg <= main_for_inc_15_storemerge_storemerge;
	end
	if (((cur_state == LEGUP_F_main_BB_NodeBlock1_25) & (fsm_stall == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge_reg <= main_for_inc_15_storemerge_storemerge;
	end
	if ((((cur_state == LEGUP_F_main_BB_NodeBlock_26) & (fsm_stall == 1'd0)) & (main_NodeBlock_Pivot == 1'd0))) begin
		main_for_inc_15_storemerge_storemerge_reg <= main_for_inc_15_storemerge_storemerge;
	end
	if ((((cur_state == LEGUP_F_main_BB_LeafBlock_27) & (fsm_stall == 1'd0)) & (main_LeafBlock_SwitchLeaf == 1'd1))) begin
		main_for_inc_15_storemerge_storemerge_reg <= main_for_inc_15_storemerge_storemerge;
	end
end
always @(*) begin
		main_for_inc_15_exitcond324 = (main_for_cond43_preheader_37_reg == 32'd18);
end
always @(*) begin
		main_for_inc_15_for_cond43_preheader_crit_edge_pre = main_entry_vla2932_out_a;
end
always @(*) begin
	main_entry_dist_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_dist_i_address_a = (main_for_cond169_preheader_arrayidx1_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_dist_i_address_a = (main_for_cond169_preheader_arrayidx1_2_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_dist_i_address_a = (main_for_cond169_preheader_arrayidx1_4_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_dist_i_address_a = (main_for_cond169_preheader_arrayidx1_6_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_dist_i_address_a = (main_for_cond169_preheader_arrayidx1_8_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_dist_i_address_a = (main_for_cond169_preheader_arrayidx1_10_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_dist_i_address_a = (main_for_cond169_preheader_arrayidx1_12_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_dist_i_address_a = (main_for_cond169_preheader_arrayidx1_14_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_77)) begin
		main_entry_dist_i_address_a = (main_for_body172_arrayidx3_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true16_i_92)) begin
		main_entry_dist_i_address_a = (main_minDistance_exit_i_arrayidx17_i_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_dist_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_77)) begin
		main_entry_dist_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_dist_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_dist_i_in_a = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_dist_i_in_a = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_dist_i_in_a = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_dist_i_in_a = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_dist_i_in_a = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_dist_i_in_a = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_dist_i_in_a = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_dist_i_in_a = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_77)) begin
		main_entry_dist_i_in_a = 32'd0;
	end
end
always @(*) begin
	main_entry_dist_i_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_dist_i_address_b = (main_for_cond169_preheader_arrayidx1_1_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_dist_i_address_b = (main_for_cond169_preheader_arrayidx1_3_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_dist_i_address_b = (main_for_cond169_preheader_arrayidx1_5_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_dist_i_address_b = (main_for_cond169_preheader_arrayidx1_7_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_dist_i_address_b = (main_for_cond169_preheader_arrayidx1_9_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_dist_i_address_b = (main_for_cond169_preheader_arrayidx1_11_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_dist_i_address_b = (main_for_cond169_preheader_arrayidx1_13_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_dist_i_address_b = (main_for_cond169_preheader_arrayidx1_15_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_i_82)) begin
		main_entry_dist_i_address_b = (main_land_lhs_true_i_i_arrayidx2_i_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true16_i_92)) begin
		main_entry_dist_i_address_b = (main_for_body11_i_arrayidx20_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_94)) begin
		main_entry_dist_i_address_b = (main_for_body11_i_arrayidx20_i_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_dist_i_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_94)) begin
		main_entry_dist_i_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_dist_i_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_dist_i_in_b = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_dist_i_in_b = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_dist_i_in_b = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_dist_i_in_b = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_dist_i_in_b = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_dist_i_in_b = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_dist_i_in_b = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_dist_i_in_b = 32'd2147483647;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_94)) begin
		main_entry_dist_i_in_b = main_land_lhs_true16_i_add_i_reg;
	end
end
always @(*) begin
	main_entry_sptSet_i_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_sptSet_i_address_a = (main_for_cond169_preheader_arrayidx2_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_sptSet_i_address_a = (main_for_cond169_preheader_arrayidx2_2_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_sptSet_i_address_a = (main_for_cond169_preheader_arrayidx2_4_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_sptSet_i_address_a = (main_for_cond169_preheader_arrayidx2_6_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_sptSet_i_address_a = (main_for_cond169_preheader_arrayidx2_8_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_sptSet_i_address_a = (main_for_cond169_preheader_arrayidx2_10_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_sptSet_i_address_a = (main_for_cond169_preheader_arrayidx2_12_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_sptSet_i_address_a = (main_for_cond169_preheader_arrayidx2_14_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body_i_i_80)) begin
		main_entry_sptSet_i_address_a = (main_for_body_i_i_arrayidx_i_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body11_i_87)) begin
		main_entry_sptSet_i_address_a = (main_for_body11_i_arrayidx12_i >>> 3'd2);
	end
end
always @(*) begin
	main_entry_sptSet_i_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_sptSet_i_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_sptSet_i_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_sptSet_i_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_sptSet_i_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_sptSet_i_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_sptSet_i_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_sptSet_i_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_sptSet_i_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_sptSet_i_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_sptSet_i_in_a = 32'd0;
	end
end
always @(*) begin
	main_entry_sptSet_i_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_sptSet_i_address_b = (main_for_cond169_preheader_arrayidx2_1_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_sptSet_i_address_b = (main_for_cond169_preheader_arrayidx2_3_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_sptSet_i_address_b = (main_for_cond169_preheader_arrayidx2_5_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_sptSet_i_address_b = (main_for_cond169_preheader_arrayidx2_7_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_sptSet_i_address_b = (main_for_cond169_preheader_arrayidx2_9_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_sptSet_i_address_b = (main_for_cond169_preheader_arrayidx2_11_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_sptSet_i_address_b = (main_for_cond169_preheader_arrayidx2_13_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_sptSet_i_address_b = (main_for_cond169_preheader_arrayidx2_15_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_85)) begin
		main_entry_sptSet_i_address_b = (main_minDistance_exit_i_arrayidx8_i >>> 3'd2);
	end
end
always @(*) begin
	main_entry_sptSet_i_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_sptSet_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_sptSet_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_sptSet_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_sptSet_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_sptSet_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_sptSet_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_sptSet_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_sptSet_i_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_85)) begin
		main_entry_sptSet_i_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_sptSet_i_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_sptSet_i_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_sptSet_i_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_71)) begin
		main_entry_sptSet_i_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_72)) begin
		main_entry_sptSet_i_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_73)) begin
		main_entry_sptSet_i_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_74)) begin
		main_entry_sptSet_i_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_75)) begin
		main_entry_sptSet_i_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body172_76)) begin
		main_entry_sptSet_i_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_minDistance_exit_i_85)) begin
		main_entry_sptSet_i_in_b = 32'd1;
	end
end
always @(*) begin
	main_entry_parent_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_parent_address_a = (main_for_body172_arrayidx_i >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_94)) begin
		main_entry_parent_address_a = (main_for_body11_i_arrayidx22_i_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_dijkstra_exit_98)) begin
		main_entry_parent_address_a = (main_dijkstra_exit_arrayidx181303 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then194_103)) begin
		main_entry_parent_address_a = (main_if_then194_arrayidx181 >>> 3'd2);
	end
end
always @(*) begin
	main_entry_parent_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_parent_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_94)) begin
		main_entry_parent_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_parent_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_70)) begin
		main_entry_parent_in_a = -32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then_i_94)) begin
		main_entry_parent_in_a = main_for_inc_i_i_min_index_1_i_i_reg;
	end
end
always @(*) begin
	main_entry_m1_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_entry_m1_address_a = (main_for_body75_scevgep44 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_46)) begin
		main_entry_m1_address_a = (main_for_body75_scevgep43_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_47)) begin
		main_entry_m1_address_a = (main_for_body75_scevgep42_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_48)) begin
		main_entry_m1_address_a = (main_for_body75_scevgep41_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_49)) begin
		main_entry_m1_address_a = (main_for_body75_scevgep40_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_50)) begin
		main_entry_m1_address_a = (main_for_body75_scevgep39_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_57)) begin
		main_entry_m1_address_a = (main_for_body75_scevgep32_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_59)) begin
		main_entry_m1_address_a = (main_for_body75_scevgep30_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_64)) begin
		main_entry_m1_address_a = (main_for_cond92_preheader_scevgep26 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_land_lhs_true_i_90)) begin
		main_entry_m1_address_a = (main_land_lhs_true_i_scevgep >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_110)) begin
		main_entry_m1_address_a = (main_for_cond92_preheader_scevgep22_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_111)) begin
		main_entry_m1_address_a = (main_for_cond92_preheader_scevgep20_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_entry_m1_address_a = (main_for_cond92_preheader_scevgep22_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_entry_m1_address_a = (main_for_cond92_preheader_scevgep20_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_115)) begin
		main_entry_m1_address_a = (main_for_inc163_us_3_scevgep14_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_116)) begin
		main_entry_m1_address_a = (main_for_inc163_us_3_scevgep16_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_117)) begin
		main_entry_m1_address_a = (main_for_inc163_us_3_scevgep17_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_118)) begin
		main_entry_m1_address_a = (main_for_inc163_us_3_scevgep18_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_m1_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_46)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_47)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_48)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_49)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_50)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_57)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_59)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_64)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_110)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_111)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_115)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_116)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_117)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_118)) begin
		main_entry_m1_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_m1_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_entry_m1_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_46)) begin
		main_entry_m1_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_47)) begin
		main_entry_m1_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_48)) begin
		main_entry_m1_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_49)) begin
		main_entry_m1_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_50)) begin
		main_entry_m1_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_57)) begin
		main_entry_m1_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_59)) begin
		main_entry_m1_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_64)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_110)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_111)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_115)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_116)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_117)) begin
		main_entry_m1_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_118)) begin
		main_entry_m1_in_a = 32'd1;
	end
end
always @(*) begin
	main_entry_m1_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body75_51)) begin
		main_entry_m1_address_b = (main_for_body75_scevgep38_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_52)) begin
		main_entry_m1_address_b = (main_for_body75_scevgep37_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_53)) begin
		main_entry_m1_address_b = (main_for_body75_scevgep36_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_54)) begin
		main_entry_m1_address_b = (main_for_body75_scevgep35_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_55)) begin
		main_entry_m1_address_b = (main_for_body75_scevgep34_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_56)) begin
		main_entry_m1_address_b = (main_for_body75_scevgep33_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_58)) begin
		main_entry_m1_address_b = (main_for_body75_scevgep31_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_60)) begin
		main_entry_m1_address_b = (main_for_body75_scevgep29_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_65)) begin
		main_entry_m1_address_b = (main_for_cond92_preheader_scevgep27_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_110)) begin
		main_entry_m1_address_b = (main_for_cond92_preheader_scevgep25_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_111)) begin
		main_entry_m1_address_b = (main_for_cond92_preheader_scevgep23_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_entry_m1_address_b = (main_for_cond92_preheader_scevgep25_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_entry_m1_address_b = (main_for_cond92_preheader_scevgep23_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_115)) begin
		main_entry_m1_address_b = (main_for_inc163_us_3_scevgep15_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_116)) begin
		main_entry_m1_address_b = (main_for_inc163_us_3_scevgep24_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_117)) begin
		main_entry_m1_address_b = (main_for_inc163_us_3_scevgep21_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_118)) begin
		main_entry_m1_address_b = (main_for_inc163_us_3_scevgep19_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_m1_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body75_51)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_52)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_53)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_54)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_55)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_56)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_58)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_60)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_65)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_110)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_111)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_115)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_116)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_117)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_118)) begin
		main_entry_m1_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_m1_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body75_51)) begin
		main_entry_m1_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_52)) begin
		main_entry_m1_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_53)) begin
		main_entry_m1_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_54)) begin
		main_entry_m1_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_55)) begin
		main_entry_m1_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_56)) begin
		main_entry_m1_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_58)) begin
		main_entry_m1_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_body75_60)) begin
		main_entry_m1_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_cond92_preheader_65)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_110)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_3_111)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_113)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_114)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_115)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_116)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_117)) begin
		main_entry_m1_in_b = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc163_us_3_118)) begin
		main_entry_m1_in_b = 32'd1;
	end
end
always @(*) begin
	main_entry_indice_e_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_entry_indice_e_address_a = (main_for_body75_arrayidx76 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end185_101)) begin
		main_entry_indice_e_address_a = (main_if_end185_arrayidx189 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then194_103)) begin
		main_entry_indice_e_address_a = (main_if_end185_arrayidx189_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_indice_e_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_entry_indice_e_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then194_103)) begin
		main_entry_indice_e_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_indice_e_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_entry_indice_e_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then194_103)) begin
		main_entry_indice_e_in_a = main_if_then194_add202;
	end
end
always @(*) begin
	main_entry_indice_s_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_entry_indice_s_address_a = (main_for_body75_arrayidx77 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_end185_101)) begin
		main_entry_indice_s_address_a = (main_if_end185_arrayidx186 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_if_then194_103)) begin
		main_entry_indice_s_address_a = (main_if_end185_arrayidx186_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_indice_s_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_entry_indice_s_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then194_103)) begin
		main_entry_indice_s_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_indice_s_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body75_45)) begin
		main_entry_indice_s_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_if_then194_103)) begin
		main_entry_indice_s_in_a = main_if_then194_add204;
	end
end
always @(*) begin
	main_entry_vla2932_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla2932_address_a = (main_entry_0 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla2932_address_a = (main_entry_4_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla2932_address_a = (main_entry_8_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla2932_address_a = (main_entry_12_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla2932_address_a = (main_entry_16_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla2932_address_a = (main_entry_20_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla2932_address_a = (main_entry_24_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla2932_address_a = (main_entry_28_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla2932_address_a = (main_entry_32_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc_15_for_cond43_preheader_crit_edge_130)) begin
		main_entry_vla2932_address_a = (main_for_cond43_preheader_scevgep49_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla2932_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla2932_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla2932_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla2932_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla2932_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla2932_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla2932_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla2932_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla2932_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla2932_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla2932_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla2932_in_a = 32'd14;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla2932_in_a = 32'd12;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla2932_in_a = 32'd10;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla2932_in_a = 32'd8;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla2932_in_a = 32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla2932_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla2932_in_a = 32'd7;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla2932_in_a = 32'd9;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla2932_in_a = 32'd13;
	end
end
always @(*) begin
	main_entry_vla2932_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla2932_address_b = (main_entry_2 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla2932_address_b = (main_entry_6_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla2932_address_b = (main_entry_10_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla2932_address_b = (main_entry_14_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla2932_address_b = (main_entry_18_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla2932_address_b = (main_entry_22_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla2932_address_b = (main_entry_26_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla2932_address_b = (main_entry_30_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla2932_address_b = (main_entry_34_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla2932_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla2932_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla2932_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla2932_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla2932_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla2932_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla2932_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla2932_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla2932_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla2932_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_vla2932_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla2932_in_b = 32'd14;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla2932_in_b = 32'd10;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla2932_in_b = 32'd8;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla2932_in_b = 32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla2932_in_b = 32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla2932_in_b = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla2932_in_b = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla2932_in_b = 32'd6;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla2932_in_b = 32'd11;
	end
end
always @(*) begin
	main_entry_vla12943_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla12943_address_a = (main_entry_1 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla12943_address_a = (main_entry_5_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla12943_address_a = (main_entry_9_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla12943_address_a = (main_entry_13_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla12943_address_a = (main_entry_17_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla12943_address_a = (main_entry_21_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla12943_address_a = (main_entry_25_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla12943_address_a = (main_entry_29_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla12943_address_a = (main_entry_33_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc67_15_for_cond58_preheader_crit_edge_124)) begin
		main_entry_vla12943_address_a = (main_for_cond58_preheader_scevgep47_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla12943_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla12943_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla12943_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla12943_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla12943_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla12943_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla12943_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla12943_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla12943_write_enable_a = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla12943_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla12943_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla12943_in_a = 32'd13;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla12943_in_a = 32'd10;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla12943_in_a = 32'd8;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla12943_in_a = 32'd7;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla12943_in_a = 32'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla12943_in_a = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla12943_in_a = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla12943_in_a = 32'd6;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla12943_in_a = 32'd11;
	end
end
always @(*) begin
	main_entry_vla12943_address_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla12943_address_b = (main_entry_3 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla12943_address_b = (main_entry_7_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla12943_address_b = (main_entry_11_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla12943_address_b = (main_entry_15_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla12943_address_b = (main_entry_19_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla12943_address_b = (main_entry_23_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla12943_address_b = (main_entry_27_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla12943_address_b = (main_entry_31_reg >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla12943_address_b = (main_entry_35_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla12943_write_enable_b = 'd0;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla12943_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla12943_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla12943_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla12943_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla12943_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla12943_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla12943_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla12943_write_enable_b = 1'd1;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla12943_write_enable_b = 1'd1;
	end
end
always @(*) begin
	main_entry_vla12943_in_b = 'dx;
	if ((cur_state == LEGUP_F_main_BB_entry_1)) begin
		main_entry_vla12943_in_b = 32'd12;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_2)) begin
		main_entry_vla12943_in_b = 32'd9;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_3)) begin
		main_entry_vla12943_in_b = 32'd5;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_4)) begin
		main_entry_vla12943_in_b = 32'd3;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_5)) begin
		main_entry_vla12943_in_b = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_6)) begin
		main_entry_vla12943_in_b = 32'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_7)) begin
		main_entry_vla12943_in_b = 32'd2;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_8)) begin
		main_entry_vla12943_in_b = 32'd4;
	end
	if ((cur_state == LEGUP_F_main_BB_entry_9)) begin
		main_entry_vla12943_in_b = 32'd9;
	end
end
always @(*) begin
	main_entry_vla39295_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_vla39295_address_a = (main_for_body172_arrayidx173 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc_15_storemerge_126)) begin
		main_entry_vla39295_address_a = (main_for_cond43_preheader_arrayidx49_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla39295_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_inc_15_storemerge_126)) begin
		main_entry_vla39295_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla39295_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_inc_15_storemerge_126)) begin
		main_entry_vla39295_in_a = {28'd0,main_for_inc_15_storemerge_storemerge_reg};
	end
end
always @(*) begin
	main_entry_vla40296_address_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_body172_69)) begin
		main_entry_vla40296_address_a = (main_for_body172_arrayidx174 >>> 3'd2);
	end
	if ((cur_state == LEGUP_F_main_BB_for_inc67_15_storemerge_120)) begin
		main_entry_vla40296_address_a = (main_for_cond58_preheader_arrayidx65_reg >>> 3'd2);
	end
end
always @(*) begin
	main_entry_vla40296_write_enable_a = 'd0;
	if ((cur_state == LEGUP_F_main_BB_for_inc67_15_storemerge_120)) begin
		main_entry_vla40296_write_enable_a = 1'd1;
	end
end
always @(*) begin
	main_entry_vla40296_in_a = 'dx;
	if ((cur_state == LEGUP_F_main_BB_for_inc67_15_storemerge_120)) begin
		main_entry_vla40296_in_a = {28'd0,main_for_inc67_15_storemerge_storemerge52_reg};
	end
end
assign main_for_cond43_preheader_Pivot30_op1_temp = 32'd8;
assign main_NodeBlock27_Pivot28_op1_temp = 32'd12;
assign main_NodeBlock25_Pivot26_op1_temp = 32'd14;
assign main_NodeBlock23_Pivot24_op1_temp = 32'd15;
assign main_NodeBlock19_Pivot20_op1_temp = 32'd13;
assign main_NodeBlock17_Pivot18_op1_temp = 32'd10;
assign main_NodeBlock15_Pivot16_op1_temp = 32'd11;
assign main_NodeBlock13_Pivot14_op1_temp = 32'd9;
assign main_NodeBlock11_Pivot12_op1_temp = 32'd4;
assign main_NodeBlock9_Pivot10_op1_temp = 32'd6;
assign main_NodeBlock7_Pivot8_op1_temp = 32'd7;
assign main_NodeBlock5_Pivot6_op1_temp = 32'd5;
assign main_NodeBlock3_Pivot4_op1_temp = 32'd2;
assign main_NodeBlock1_Pivot2_op1_temp = 32'd3;
assign main_NodeBlock_Pivot_op1_temp = 32'd1;
assign main_for_cond58_preheader_Pivot65_op1_temp = 32'd8;
assign main_NodeBlock62_Pivot63_op1_temp = 32'd12;
assign main_NodeBlock60_Pivot61_op1_temp = 32'd14;
assign main_NodeBlock58_Pivot59_op1_temp = 32'd15;
assign main_NodeBlock54_Pivot55_op1_temp = 32'd13;
assign main_NodeBlock52_Pivot53_op1_temp = 32'd10;
assign main_NodeBlock50_Pivot51_op1_temp = 32'd11;
assign main_NodeBlock48_Pivot49_op1_temp = 32'd9;
assign main_NodeBlock46_Pivot47_op1_temp = 32'd4;
assign main_NodeBlock44_Pivot45_op1_temp = 32'd6;
assign main_NodeBlock42_Pivot43_op1_temp = 32'd7;
assign main_NodeBlock40_Pivot41_op1_temp = 32'd5;
assign main_NodeBlock38_Pivot39_op1_temp = 32'd2;
assign main_NodeBlock36_Pivot37_op1_temp = 32'd3;
assign main_NodeBlock34_Pivot35_op1_temp = 32'd1;
always @(*) begin
	main_for_body75_i_0312_reg_width_extended = {23'd0,main_for_body75_i_0312_reg};
end
assign main_for_body75_bit_concat23_bit_select_operand_2 = 4'd0;
assign main_for_body75_bit_concat22_bit_select_operand_2 = 4'd1;
assign main_for_body75_bit_concat21_bit_select_operand_2 = 4'd2;
assign main_for_body75_bit_concat20_bit_select_operand_2 = 4'd3;
assign main_for_body75_bit_concat19_bit_select_operand_2 = 4'd4;
assign main_for_body75_bit_concat18_bit_select_operand_2 = 4'd5;
assign main_for_body75_bit_concat17_bit_select_operand_2 = 4'd6;
assign main_for_body75_bit_concat16_bit_select_operand_2 = 4'd7;
assign main_for_body75_bit_concat15_bit_select_operand_2 = -4'd8;
assign main_for_body75_bit_concat14_bit_select_operand_2 = -4'd7;
assign main_for_body75_bit_concat13_bit_select_operand_2 = -4'd6;
assign main_for_body75_bit_concat12_bit_select_operand_2 = -4'd5;
assign main_for_body75_bit_concat11_bit_select_operand_2 = -4'd4;
assign main_for_body75_bit_concat10_bit_select_operand_2 = -4'd3;
assign main_for_body75_bit_concat9_bit_select_operand_2 = -4'd2;
assign main_for_body75_bit_concat8_bit_select_operand_2 = -4'd1;
always @(*) begin
	main_for_cond92_preheader_43_reg_width_extended = {27'd0,main_for_cond92_preheader_43_reg};
end
assign main_for_cond92_preheader_bit_concat6_bit_select_operand_2 = 2'd0;
assign main_for_cond92_preheader_bit_concat4_bit_select_operand_2 = 6'd0;
assign main_for_cond92_preheader_bit_concat2_bit_select_operand_2 = 1'd1;
always @(*) begin
	main_for_cond92_preheader_cmp95_op0_temp = {1'd0,main_for_cond92_preheader_43_reg};
end
assign main_for_cond92_preheader_cmp95_op1_temp = 32'd3;
assign main_minDistance_exit_i_bit_concat_bit_select_operand_2 = 4'd0;
assign main_if_end185_cmp187_op1_temp = 32'd4;
assign main_if_end185_cmp190_op1_temp = 32'd4;
always @(*) begin
	main_for_inc212_cmp170_op0_temp = {1'd0,main_for_body172_inc213_reg};
end
assign main_for_inc212_cmp170_op1_temp = 32'd19;
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		finish <= 1'd0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end214_109)) begin
		finish <= (fsm_stall == 1'd0);
	end
end
always @(posedge clk) begin
	if ((cur_state == LEGUP_0)) begin
		return_val <= 0;
	end
	if ((cur_state == LEGUP_F_main_BB_for_end214_109)) begin
		return_val <= 32'd0;
	end
end

endmodule
module ram_dual_port
(
	clk,
	clken,
	address_a,
	address_b,
	wren_a,
	data_a,
	byteena_a,
	wren_b,
	data_b,
	byteena_b,
	q_b,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  width_b = 1'd0;
parameter  widthad_b = 1'd0;
parameter  numwords_b = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
parameter  width_be_b = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input [(widthad_b-1):0] address_b;
output wire [(width_b-1):0] q_b;
wire [(width_b-1):0] q_b_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
input  wren_b;
input [(width_b-1):0] data_b;
input [width_be_b-1:0] byteena_b;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
	.address_b (address_b),
    .addressstall_b (1'd0),
    .rden_b (clken),
    .q_b (q_b),
    .wren_a (wren_a),
    .data_a (data_a),
    .wren_b (wren_b),
    .data_b (data_b),
    .byteena_b (byteena_b),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.width_byteena_b = width_be_b,
    altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "Arria10",
    altsyncram_component.clock_enable_input_b = "BYPASS",
    altsyncram_component.clock_enable_output_b = "BYPASS",
    altsyncram_component.outdata_aclr_b = "NONE",
    altsyncram_component.outdata_reg_b = output_registered,
    altsyncram_component.numwords_b = numwords_b,
    altsyncram_component.widthad_b = widthad_b,
    altsyncram_component.width_b = width_b,
    altsyncram_component.address_reg_b = "CLOCK0",
    altsyncram_component.byteena_reg_b = "CLOCK0",
    altsyncram_component.indata_reg_b = "CLOCK0",
    altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
module ram_single_port_intel
(
	clk,
	clken,
	address_a,
	wren_a,
	data_a,
	byteena_a,
	q_a
);

parameter  width_a = 1'd0;
parameter  widthad_a = 1'd0;
parameter  numwords_a = 1'd0;
parameter  latency = 1;
parameter  init_file = "UNUSED";
parameter  width_be_a = 1'd0;
localparam output_registered = (latency == 1)? "UNREGISTERED" : "CLOCK0";
input  clk;
input  clken;
input [(widthad_a-1):0] address_a;
output wire [(width_a-1):0] q_a;
wire [(width_a-1):0] q_a_wire;
input  wren_a;
input [(width_a-1):0] data_a;
input [width_be_a-1:0] byteena_a;
reg  clk_wire;

altsyncram altsyncram_component (
	.address_a (address_a),
    .clock0 (clk_wire),
    .clock1 (1'd1),
    .clocken0 (clken),
    .clocken1 (1'd1),
    .clocken2 (1'd1),
    .clocken3 (1'd1),
    .aclr0 (1'd0),
    .aclr1 (1'd0),
    .addressstall_a (1'd0),
    .eccstatus (),
    .rden_a (clken),
    .q_a (q_a),
    .wren_a (wren_a),
    .data_a (data_a),
    .byteena_a (byteena_a)
);
defparam
    altsyncram_component.width_byteena_a = width_be_a,
    altsyncram_component.operation_mode = "SINGLE_PORT",
    altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
    altsyncram_component.init_file = init_file,
    altsyncram_component.lpm_hint = "ENABLE_RUNTIME_MOD=NO",
    altsyncram_component.lpm_type = "altsyncram",
    altsyncram_component.power_up_uninitialized = "FALSE",
    altsyncram_component.intended_device_family = "Arria10",
    altsyncram_component.clock_enable_input_a = "BYPASS",
    altsyncram_component.clock_enable_output_a = "BYPASS",
    altsyncram_component.outdata_aclr_a = "NONE",
    altsyncram_component.outdata_reg_a = output_registered,
    altsyncram_component.numwords_a = numwords_a,
    altsyncram_component.widthad_a = widthad_a,
    altsyncram_component.width_a = width_a;

always @(*) begin
	clk_wire = clk;
end


endmodule
`timescale 1 ns / 1 ns
module main_tb
(
);

reg  clk;
reg  reset;
reg  start;
wire [31:0] return_val;
wire  finish;


top top_inst (
	.clk (clk),
	.reset (reset),
	.start (start),
	.finish (finish),
	.return_val (return_val)
);




initial 
    clk = 0;
always @(clk)
    clk <= #10 ~clk;

initial begin
//$monitor("At t=%t clk=%b %b %b %b %d", $time, clk, reset, start, finish, return_val);
reset <= 1;
@(negedge clk);
reset <= 0;
start <= 1;
@(negedge clk);
start <= 0;
end

always@(posedge clk) begin
    if (finish == 1) begin
        $display("At t=%t clk=%b finish=%b return_val=%d", $time, clk, finish, return_val);
        $display("Cycles: %d", ($time-50)/20);
        $finish;
    end
end


endmodule
